module polar_decoder (
    clk,
    rst_n,
    module_en,
    proc_done,
    raddr,
    rdata,
    waddr,
    wdata
);
// IO description
input  wire         clk;
input  wire         rst_n;
input  wire         module_en;
input  wire [191:0] rdata;
output wire [ 10:0] raddr;
output wire [  5:0] waddr;
output wire [139:0] wdata;
output wire         proc_done;

// **************************//
// *****   DECLARATION  *****//
// **************************//

reg         en;
reg [191:0] in_data;

reg       firstRead;
reg [5:0] n_package;
reg [9:0] N;
reg [7:0] K;

reg [2:0] state, state_nxt;
reg [9:0] counter;
reg [5:0] counter_p;
parameter IDLE	 = 3'd0;
parameter SUB 	 = 3'd1;
parameter SUB2   = 3'd2;
parameter READ	 = 3'd3;
parameter DECODE = 3'd4;
parameter DONE	 = 3'd5;

integer i;

parameter LLR_bit = 18;
reg [(LLR_bit-1):0] LLR [512:1];

reg  [511:0] frozen;
reg    [1:0] usum2;
reg    [3:0] usum4;
reg    [7:0] usum8;
reg   [15:0] usum16;
reg   [31:0] usum32;
reg   [63:0] usum64;
reg  [127:0] usum128;
reg  [255:0] usum256;
reg  [255:0] u;
reg  [139:0] answer;

wire [10:0] u_counter = (counter>>1);
wire [10:0] usum_counter = counter - (counter>>1);
wire [10:0] usum_counter_minus = counter - (counter>>1) - 1;

wire [255:0] usum_256;
wire [127:0] usum_128;
wire  [63:0] usum_64;
wire  [31:0] usum_32;
wire  [15:0] usum_16;
wire   [7:0] usum_8;
wire   [3:0] usum_4;
wire   [1:0] usum_2;

wire signed [(LLR_bit-1):0] input1_128;
wire signed [(LLR_bit-1):0] input2_128;
wire signed [(LLR_bit-1):0] input1_256;
wire signed [(LLR_bit-1):0] input2_256;
wire signed [(LLR_bit-1):0] input1_512;
wire signed [(LLR_bit-1):0] input2_512;

wire [1:0] pnode_128;
wire [1:0] pnode_256;
wire [1:0] pnode_512;
wire [1:0] pnode_N;

reg [7:0] counter_answer;

reg   [5:0] waddr_r;
reg [139:0] wdata_r;
reg         proc_done_r;

// *******************//
// *****   FSM   *****//
// *******************//

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        en      <= 0;
        in_data <= 0;
    end else if(proc_done_r) begin
        en      <= 0;
        in_data <= 0;
    end else begin
        en      <= module_en;
        in_data <= rdata;
    end
end

always @(*) begin
    case(state)
        IDLE:    state_nxt = (en) ? SUB : IDLE;
        SUB:	 state_nxt = SUB2;
        SUB2:	 state_nxt = READ;
        READ:    state_nxt = (counter == 33) ? DECODE: READ;
        DECODE:  state_nxt = (counter == N-1) ? DONE : DECODE;
        DONE:    state_nxt = SUB;
		default: state_nxt = IDLE;
    endcase
end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        state     <= IDLE;
        firstRead <= 1;
        n_package <= 0;
        N         <= 0;
        K         <= 0;
        counter   <= 0;
        counter_p <= 0;
    end else if(proc_done_r) begin
        state     <= IDLE;
        firstRead <= 1;
        n_package <= 0;
        N         <= 0;
        K         <= 0;
        counter   <= 0;
        counter_p <= 0;
    end else begin
        state     <= state_nxt;
        firstRead <= (state == READ) ? 0 : firstRead;
        n_package <= (state == READ && counter == 0 && firstRead) ? in_data[6:0] : n_package;
        N         <= (state == READ && counter == 1) ? in_data[9:0] : N;
        K         <= (state == READ && counter == 1) ? in_data[17:10] : K;
        counter   <= (state == state_nxt) ? counter+1 : 0;
        counter_p <= (state == DONE) ? counter_p+1 : counter_p;
    end
end

// ***********************//
// **** PREPROCESSING ****//
// ***********************//

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		for(i=1; i<=512; i=i+1)
			LLR[i] <= 0;
	end else if (state==READ && 2<=counter && counter<=33) begin
		case (counter) // synopsys full_case
			2:  begin for(i=1; i<=16; i=i+1) LLR[i]     <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			3:  begin for(i=1; i<=16; i=i+1) LLR[i+16]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			4:  begin for(i=1; i<=16; i=i+1) LLR[i+32]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			5:  begin for(i=1; i<=16; i=i+1) LLR[i+48]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			6:  begin for(i=1; i<=16; i=i+1) LLR[i+64]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			7:  begin for(i=1; i<=16; i=i+1) LLR[i+80]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			8:  begin for(i=1; i<=16; i=i+1) LLR[i+96]  <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			9:  begin for(i=1; i<=16; i=i+1) LLR[i+112] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			10: begin for(i=1; i<=16; i=i+1) LLR[i+128] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			11: begin for(i=1; i<=16; i=i+1) LLR[i+144] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			12: begin for(i=1; i<=16; i=i+1) LLR[i+160] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			13: begin for(i=1; i<=16; i=i+1) LLR[i+176] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			14: begin for(i=1; i<=16; i=i+1) LLR[i+192] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			15: begin for(i=1; i<=16; i=i+1) LLR[i+208] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			16: begin for(i=1; i<=16; i=i+1) LLR[i+224] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			17: begin for(i=1; i<=16; i=i+1) LLR[i+240] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			18: begin for(i=1; i<=16; i=i+1) LLR[i+256] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			19: begin for(i=1; i<=16; i=i+1) LLR[i+272] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			20: begin for(i=1; i<=16; i=i+1) LLR[i+288] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			21: begin for(i=1; i<=16; i=i+1) LLR[i+304] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			22: begin for(i=1; i<=16; i=i+1) LLR[i+320] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			23: begin for(i=1; i<=16; i=i+1) LLR[i+336] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			24: begin for(i=1; i<=16; i=i+1) LLR[i+352] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			25: begin for(i=1; i<=16; i=i+1) LLR[i+368] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			26: begin for(i=1; i<=16; i=i+1) LLR[i+384] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			27: begin for(i=1; i<=16; i=i+1) LLR[i+400] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			28: begin for(i=1; i<=16; i=i+1) LLR[i+416] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			29: begin for(i=1; i<=16; i=i+1) LLR[i+432] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			30: begin for(i=1; i<=16; i=i+1) LLR[i+448] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			31: begin for(i=1; i<=16; i=i+1) LLR[i+464] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			32: begin for(i=1; i<=16; i=i+1) LLR[i+480] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
			33: begin for(i=1; i<=16; i=i+1) LLR[i+496] <={{(LLR_bit-12){in_data[(i*12-1)]}}, in_data[(i*12-1) -: 12]}; end
		endcase
	end else begin
		for(i=1; i<=512; i=i+1)
			LLR[i] <= LLR[i];
	end
end

// ***********************//
// *****   DECODER   *****//
// ***********************//

assign usum_256 = {u[255],u[255]^u[127],u[255]^u[191],u[255]^u[191]^u[127]^u[63],u[255]^u[223],u[255]^u[223]^u[127]^u[95],u[255]^u[223]^u[191]^u[159],u[255]^u[223]^u[191]^u[159]^u[127]^u[95]^u[63]^u[31],u[255]^u[239],u[255]^u[239]^u[127]^u[111],u[255]^u[239]^u[191]^u[175],u[255]^u[239]^u[191]^u[175]^u[127]^u[111]^u[63]^u[47],u[255]^u[239]^u[223]^u[207],u[255]^u[239]^u[223]^u[207]^u[127]^u[111]^u[95]^u[79],u[255]^u[239]^u[223]^u[207]^u[191]^u[175]^u[159]^u[143],u[255]^u[239]^u[223]^u[207]^u[191]^u[175]^u[159]^u[143]^u[127]^u[111]^u[95]^u[79]^u[63]^u[47]^u[31]^u[15],u[255]^u[247],u[255]^u[247]^u[127]^u[119],u[255]^u[247]^u[191]^u[183],u[255]^u[247]^u[191]^u[183]^u[127]^u[119]^u[63]^u[55],u[255]^u[247]^u[223]^u[215],u[255]^u[247]^u[223]^u[215]^u[127]^u[119]^u[95]^u[87],u[255]^u[247]^u[223]^u[215]^u[191]^u[183]^u[159]^u[151],u[255]^u[247]^u[223]^u[215]^u[191]^u[183]^u[159]^u[151]^u[127]^u[119]^u[95]^u[87]^u[63]^u[55]^u[31]^u[23],u[255]^u[247]^u[239]^u[231],u[255]^u[247]^u[239]^u[231]^u[127]^u[119]^u[111]^u[103],u[255]^u[247]^u[239]^u[231]^u[191]^u[183]^u[175]^u[167],u[255]^u[247]^u[239]^u[231]^u[191]^u[183]^u[175]^u[167]^u[127]^u[119]^u[111]^u[103]^u[63]^u[55]^u[47]^u[39],u[255]^u[247]^u[239]^u[231]^u[223]^u[215]^u[207]^u[199],u[255]^u[247]^u[239]^u[231]^u[223]^u[215]^u[207]^u[199]^u[127]^u[119]^u[111]^u[103]^u[95]^u[87]^u[79]^u[71],u[255]^u[247]^u[239]^u[231]^u[223]^u[215]^u[207]^u[199]^u[191]^u[183]^u[175]^u[167]^u[159]^u[151]^u[143]^u[135],u[255]^u[247]^u[239]^u[231]^u[223]^u[215]^u[207]^u[199]^u[191]^u[183]^u[175]^u[167]^u[159]^u[151]^u[143]^u[135]^u[127]^u[119]^u[111]^u[103]^u[95]^u[87]^u[79]^u[71]^u[63]^u[55]^u[47]^u[39]^u[31]^u[23]^u[15]^u[7],u[255]^u[251],u[255]^u[251]^u[127]^u[123],u[255]^u[251]^u[191]^u[187],u[255]^u[251]^u[191]^u[187]^u[127]^u[123]^u[63]^u[59],u[255]^u[251]^u[223]^u[219],u[255]^u[251]^u[223]^u[219]^u[127]^u[123]^u[95]^u[91],u[255]^u[251]^u[223]^u[219]^u[191]^u[187]^u[159]^u[155],u[255]^u[251]^u[223]^u[219]^u[191]^u[187]^u[159]^u[155]^u[127]^u[123]^u[95]^u[91]^u[63]^u[59]^u[31]^u[27],u[255]^u[251]^u[239]^u[235],u[255]^u[251]^u[239]^u[235]^u[127]^u[123]^u[111]^u[107],u[255]^u[251]^u[239]^u[235]^u[191]^u[187]^u[175]^u[171],u[255]^u[251]^u[239]^u[235]^u[191]^u[187]^u[175]^u[171]^u[127]^u[123]^u[111]^u[107]^u[63]^u[59]^u[47]^u[43],u[255]^u[251]^u[239]^u[235]^u[223]^u[219]^u[207]^u[203],u[255]^u[251]^u[239]^u[235]^u[223]^u[219]^u[207]^u[203]^u[127]^u[123]^u[111]^u[107]^u[95]^u[91]^u[79]^u[75],u[255]^u[251]^u[239]^u[235]^u[223]^u[219]^u[207]^u[203]^u[191]^u[187]^u[175]^u[171]^u[159]^u[155]^u[143]^u[139],u[255]^u[251]^u[239]^u[235]^u[223]^u[219]^u[207]^u[203]^u[191]^u[187]^u[175]^u[171]^u[159]^u[155]^u[143]^u[139]^u[127]^u[123]^u[111]^u[107]^u[95]^u[91]^u[79]^u[75]^u[63]^u[59]^u[47]^u[43]^u[31]^u[27]^u[15]^u[11],u[255]^u[251]^u[247]^u[243],u[255]^u[251]^u[247]^u[243]^u[127]^u[123]^u[119]^u[115],u[255]^u[251]^u[247]^u[243]^u[191]^u[187]^u[183]^u[179],u[255]^u[251]^u[247]^u[243]^u[191]^u[187]^u[183]^u[179]^u[127]^u[123]^u[119]^u[115]^u[63]^u[59]^u[55]^u[51],u[255]^u[251]^u[247]^u[243]^u[223]^u[219]^u[215]^u[211],u[255]^u[251]^u[247]^u[243]^u[223]^u[219]^u[215]^u[211]^u[127]^u[123]^u[119]^u[115]^u[95]^u[91]^u[87]^u[83],u[255]^u[251]^u[247]^u[243]^u[223]^u[219]^u[215]^u[211]^u[191]^u[187]^u[183]^u[179]^u[159]^u[155]^u[151]^u[147],u[255]^u[251]^u[247]^u[243]^u[223]^u[219]^u[215]^u[211]^u[191]^u[187]^u[183]^u[179]^u[159]^u[155]^u[151]^u[147]^u[127]^u[123]^u[119]^u[115]^u[95]^u[91]^u[87]^u[83]^u[63]^u[59]^u[55]^u[51]^u[31]^u[27]^u[23]^u[19],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[127]^u[123]^u[119]^u[115]^u[111]^u[107]^u[103]^u[99],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[191]^u[187]^u[183]^u[179]^u[175]^u[171]^u[167]^u[163],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[191]^u[187]^u[183]^u[179]^u[175]^u[171]^u[167]^u[163]^u[127]^u[123]^u[119]^u[115]^u[111]^u[107]^u[103]^u[99]^u[63]^u[59]^u[55]^u[51]^u[47]^u[43]^u[39]^u[35],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[223]^u[219]^u[215]^u[211]^u[207]^u[203]^u[199]^u[195],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[223]^u[219]^u[215]^u[211]^u[207]^u[203]^u[199]^u[195]^u[127]^u[123]^u[119]^u[115]^u[111]^u[107]^u[103]^u[99]^u[95]^u[91]^u[87]^u[83]^u[79]^u[75]^u[71]^u[67],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[223]^u[219]^u[215]^u[211]^u[207]^u[203]^u[199]^u[195]^u[191]^u[187]^u[183]^u[179]^u[175]^u[171]^u[167]^u[163]^u[159]^u[155]^u[151]^u[147]^u[143]^u[139]^u[135]^u[131],u[255]^u[251]^u[247]^u[243]^u[239]^u[235]^u[231]^u[227]^u[223]^u[219]^u[215]^u[211]^u[207]^u[203]^u[199]^u[195]^u[191]^u[187]^u[183]^u[179]^u[175]^u[171]^u[167]^u[163]^u[159]^u[155]^u[151]^u[147]^u[143]^u[139]^u[135]^u[131]^u[127]^u[123]^u[119]^u[115]^u[111]^u[107]^u[103]^u[99]^u[95]^u[91]^u[87]^u[83]^u[79]^u[75]^u[71]^u[67]^u[63]^u[59]^u[55]^u[51]^u[47]^u[43]^u[39]^u[35]^u[31]^u[27]^u[23]^u[19]^u[15]^u[11]^u[7]^u[3],u[255]^u[253],u[255]^u[253]^u[127]^u[125],u[255]^u[253]^u[191]^u[189],u[255]^u[253]^u[191]^u[189]^u[127]^u[125]^u[63]^u[61],u[255]^u[253]^u[223]^u[221],u[255]^u[253]^u[223]^u[221]^u[127]^u[125]^u[95]^u[93],u[255]^u[253]^u[223]^u[221]^u[191]^u[189]^u[159]^u[157],u[255]^u[253]^u[223]^u[221]^u[191]^u[189]^u[159]^u[157]^u[127]^u[125]^u[95]^u[93]^u[63]^u[61]^u[31]^u[29],u[255]^u[253]^u[239]^u[237],u[255]^u[253]^u[239]^u[237]^u[127]^u[125]^u[111]^u[109],u[255]^u[253]^u[239]^u[237]^u[191]^u[189]^u[175]^u[173],u[255]^u[253]^u[239]^u[237]^u[191]^u[189]^u[175]^u[173]^u[127]^u[125]^u[111]^u[109]^u[63]^u[61]^u[47]^u[45],u[255]^u[253]^u[239]^u[237]^u[223]^u[221]^u[207]^u[205],u[255]^u[253]^u[239]^u[237]^u[223]^u[221]^u[207]^u[205]^u[127]^u[125]^u[111]^u[109]^u[95]^u[93]^u[79]^u[77],u[255]^u[253]^u[239]^u[237]^u[223]^u[221]^u[207]^u[205]^u[191]^u[189]^u[175]^u[173]^u[159]^u[157]^u[143]^u[141],u[255]^u[253]^u[239]^u[237]^u[223]^u[221]^u[207]^u[205]^u[191]^u[189]^u[175]^u[173]^u[159]^u[157]^u[143]^u[141]^u[127]^u[125]^u[111]^u[109]^u[95]^u[93]^u[79]^u[77]^u[63]^u[61]^u[47]^u[45]^u[31]^u[29]^u[15]^u[13],u[255]^u[253]^u[247]^u[245],u[255]^u[253]^u[247]^u[245]^u[127]^u[125]^u[119]^u[117],u[255]^u[253]^u[247]^u[245]^u[191]^u[189]^u[183]^u[181],u[255]^u[253]^u[247]^u[245]^u[191]^u[189]^u[183]^u[181]^u[127]^u[125]^u[119]^u[117]^u[63]^u[61]^u[55]^u[53],u[255]^u[253]^u[247]^u[245]^u[223]^u[221]^u[215]^u[213],u[255]^u[253]^u[247]^u[245]^u[223]^u[221]^u[215]^u[213]^u[127]^u[125]^u[119]^u[117]^u[95]^u[93]^u[87]^u[85],u[255]^u[253]^u[247]^u[245]^u[223]^u[221]^u[215]^u[213]^u[191]^u[189]^u[183]^u[181]^u[159]^u[157]^u[151]^u[149],u[255]^u[253]^u[247]^u[245]^u[223]^u[221]^u[215]^u[213]^u[191]^u[189]^u[183]^u[181]^u[159]^u[157]^u[151]^u[149]^u[127]^u[125]^u[119]^u[117]^u[95]^u[93]^u[87]^u[85]^u[63]^u[61]^u[55]^u[53]^u[31]^u[29]^u[23]^u[21],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[127]^u[125]^u[119]^u[117]^u[111]^u[109]^u[103]^u[101],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[191]^u[189]^u[183]^u[181]^u[175]^u[173]^u[167]^u[165],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[191]^u[189]^u[183]^u[181]^u[175]^u[173]^u[167]^u[165]^u[127]^u[125]^u[119]^u[117]^u[111]^u[109]^u[103]^u[101]^u[63]^u[61]^u[55]^u[53]^u[47]^u[45]^u[39]^u[37],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[223]^u[221]^u[215]^u[213]^u[207]^u[205]^u[199]^u[197],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[223]^u[221]^u[215]^u[213]^u[207]^u[205]^u[199]^u[197]^u[127]^u[125]^u[119]^u[117]^u[111]^u[109]^u[103]^u[101]^u[95]^u[93]^u[87]^u[85]^u[79]^u[77]^u[71]^u[69],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[223]^u[221]^u[215]^u[213]^u[207]^u[205]^u[199]^u[197]^u[191]^u[189]^u[183]^u[181]^u[175]^u[173]^u[167]^u[165]^u[159]^u[157]^u[151]^u[149]^u[143]^u[141]^u[135]^u[133],u[255]^u[253]^u[247]^u[245]^u[239]^u[237]^u[231]^u[229]^u[223]^u[221]^u[215]^u[213]^u[207]^u[205]^u[199]^u[197]^u[191]^u[189]^u[183]^u[181]^u[175]^u[173]^u[167]^u[165]^u[159]^u[157]^u[151]^u[149]^u[143]^u[141]^u[135]^u[133]^u[127]^u[125]^u[119]^u[117]^u[111]^u[109]^u[103]^u[101]^u[95]^u[93]^u[87]^u[85]^u[79]^u[77]^u[71]^u[69]^u[63]^u[61]^u[55]^u[53]^u[47]^u[45]^u[39]^u[37]^u[31]^u[29]^u[23]^u[21]^u[15]^u[13]^u[7]^u[5],u[255]^u[253]^u[251]^u[249],u[255]^u[253]^u[251]^u[249]^u[127]^u[125]^u[123]^u[121],u[255]^u[253]^u[251]^u[249]^u[191]^u[189]^u[187]^u[185],u[255]^u[253]^u[251]^u[249]^u[191]^u[189]^u[187]^u[185]^u[127]^u[125]^u[123]^u[121]^u[63]^u[61]^u[59]^u[57],u[255]^u[253]^u[251]^u[249]^u[223]^u[221]^u[219]^u[217],u[255]^u[253]^u[251]^u[249]^u[223]^u[221]^u[219]^u[217]^u[127]^u[125]^u[123]^u[121]^u[95]^u[93]^u[91]^u[89],u[255]^u[253]^u[251]^u[249]^u[223]^u[221]^u[219]^u[217]^u[191]^u[189]^u[187]^u[185]^u[159]^u[157]^u[155]^u[153],u[255]^u[253]^u[251]^u[249]^u[223]^u[221]^u[219]^u[217]^u[191]^u[189]^u[187]^u[185]^u[159]^u[157]^u[155]^u[153]^u[127]^u[125]^u[123]^u[121]^u[95]^u[93]^u[91]^u[89]^u[63]^u[61]^u[59]^u[57]^u[31]^u[29]^u[27]^u[25],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[127]^u[125]^u[123]^u[121]^u[111]^u[109]^u[107]^u[105],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[191]^u[189]^u[187]^u[185]^u[175]^u[173]^u[171]^u[169],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[191]^u[189]^u[187]^u[185]^u[175]^u[173]^u[171]^u[169]^u[127]^u[125]^u[123]^u[121]^u[111]^u[109]^u[107]^u[105]^u[63]^u[61]^u[59]^u[57]^u[47]^u[45]^u[43]^u[41],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[223]^u[221]^u[219]^u[217]^u[207]^u[205]^u[203]^u[201],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[223]^u[221]^u[219]^u[217]^u[207]^u[205]^u[203]^u[201]^u[127]^u[125]^u[123]^u[121]^u[111]^u[109]^u[107]^u[105]^u[95]^u[93]^u[91]^u[89]^u[79]^u[77]^u[75]^u[73],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[223]^u[221]^u[219]^u[217]^u[207]^u[205]^u[203]^u[201]^u[191]^u[189]^u[187]^u[185]^u[175]^u[173]^u[171]^u[169]^u[159]^u[157]^u[155]^u[153]^u[143]^u[141]^u[139]^u[137],u[255]^u[253]^u[251]^u[249]^u[239]^u[237]^u[235]^u[233]^u[223]^u[221]^u[219]^u[217]^u[207]^u[205]^u[203]^u[201]^u[191]^u[189]^u[187]^u[185]^u[175]^u[173]^u[171]^u[169]^u[159]^u[157]^u[155]^u[153]^u[143]^u[141]^u[139]^u[137]^u[127]^u[125]^u[123]^u[121]^u[111]^u[109]^u[107]^u[105]^u[95]^u[93]^u[91]^u[89]^u[79]^u[77]^u[75]^u[73]^u[63]^u[61]^u[59]^u[57]^u[47]^u[45]^u[43]^u[41]^u[31]^u[29]^u[27]^u[25]^u[15]^u[13]^u[11]^u[9],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[63]^u[61]^u[59]^u[57]^u[55]^u[53]^u[51]^u[49],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[95]^u[93]^u[91]^u[89]^u[87]^u[85]^u[83]^u[81],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[159]^u[157]^u[155]^u[153]^u[151]^u[149]^u[147]^u[145],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[159]^u[157]^u[155]^u[153]^u[151]^u[149]^u[147]^u[145]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[95]^u[93]^u[91]^u[89]^u[87]^u[85]^u[83]^u[81]^u[63]^u[61]^u[59]^u[57]^u[55]^u[53]^u[51]^u[49]^u[31]^u[29]^u[27]^u[25]^u[23]^u[21]^u[19]^u[17],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[111]^u[109]^u[107]^u[105]^u[103]^u[101]^u[99]^u[97],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[175]^u[173]^u[171]^u[169]^u[167]^u[165]^u[163]^u[161],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[175]^u[173]^u[171]^u[169]^u[167]^u[165]^u[163]^u[161]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[111]^u[109]^u[107]^u[105]^u[103]^u[101]^u[99]^u[97]^u[63]^u[61]^u[59]^u[57]^u[55]^u[53]^u[51]^u[49]^u[47]^u[45]^u[43]^u[41]^u[39]^u[37]^u[35]^u[33],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[207]^u[205]^u[203]^u[201]^u[199]^u[197]^u[195]^u[193],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[207]^u[205]^u[203]^u[201]^u[199]^u[197]^u[195]^u[193]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[111]^u[109]^u[107]^u[105]^u[103]^u[101]^u[99]^u[97]^u[95]^u[93]^u[91]^u[89]^u[87]^u[85]^u[83]^u[81]^u[79]^u[77]^u[75]^u[73]^u[71]^u[69]^u[67]^u[65],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[207]^u[205]^u[203]^u[201]^u[199]^u[197]^u[195]^u[193]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[175]^u[173]^u[171]^u[169]^u[167]^u[165]^u[163]^u[161]^u[159]^u[157]^u[155]^u[153]^u[151]^u[149]^u[147]^u[145]^u[143]^u[141]^u[139]^u[137]^u[135]^u[133]^u[131]^u[129],u[255]^u[253]^u[251]^u[249]^u[247]^u[245]^u[243]^u[241]^u[239]^u[237]^u[235]^u[233]^u[231]^u[229]^u[227]^u[225]^u[223]^u[221]^u[219]^u[217]^u[215]^u[213]^u[211]^u[209]^u[207]^u[205]^u[203]^u[201]^u[199]^u[197]^u[195]^u[193]^u[191]^u[189]^u[187]^u[185]^u[183]^u[181]^u[179]^u[177]^u[175]^u[173]^u[171]^u[169]^u[167]^u[165]^u[163]^u[161]^u[159]^u[157]^u[155]^u[153]^u[151]^u[149]^u[147]^u[145]^u[143]^u[141]^u[139]^u[137]^u[135]^u[133]^u[131]^u[129]^u[127]^u[125]^u[123]^u[121]^u[119]^u[117]^u[115]^u[113]^u[111]^u[109]^u[107]^u[105]^u[103]^u[101]^u[99]^u[97]^u[95]^u[93]^u[91]^u[89]^u[87]^u[85]^u[83]^u[81]^u[79]^u[77]^u[75]^u[73]^u[71]^u[69]^u[67]^u[65]^u[63]^u[61]^u[59]^u[57]^u[55]^u[53]^u[51]^u[49]^u[47]^u[45]^u[43]^u[41]^u[39]^u[37]^u[35]^u[33]^u[31]^u[29]^u[27]^u[25]^u[23]^u[21]^u[19]^u[17]^u[15]^u[13]^u[11]^u[9]^u[7]^u[5]^u[3]^u[1],u[255]^u[254],u[255]^u[254]^u[127]^u[126],u[255]^u[254]^u[191]^u[190],u[255]^u[254]^u[191]^u[190]^u[127]^u[126]^u[63]^u[62],u[255]^u[254]^u[223]^u[222],u[255]^u[254]^u[223]^u[222]^u[127]^u[126]^u[95]^u[94],u[255]^u[254]^u[223]^u[222]^u[191]^u[190]^u[159]^u[158],u[255]^u[254]^u[223]^u[222]^u[191]^u[190]^u[159]^u[158]^u[127]^u[126]^u[95]^u[94]^u[63]^u[62]^u[31]^u[30],u[255]^u[254]^u[239]^u[238],u[255]^u[254]^u[239]^u[238]^u[127]^u[126]^u[111]^u[110],u[255]^u[254]^u[239]^u[238]^u[191]^u[190]^u[175]^u[174],u[255]^u[254]^u[239]^u[238]^u[191]^u[190]^u[175]^u[174]^u[127]^u[126]^u[111]^u[110]^u[63]^u[62]^u[47]^u[46],u[255]^u[254]^u[239]^u[238]^u[223]^u[222]^u[207]^u[206],u[255]^u[254]^u[239]^u[238]^u[223]^u[222]^u[207]^u[206]^u[127]^u[126]^u[111]^u[110]^u[95]^u[94]^u[79]^u[78],u[255]^u[254]^u[239]^u[238]^u[223]^u[222]^u[207]^u[206]^u[191]^u[190]^u[175]^u[174]^u[159]^u[158]^u[143]^u[142],u[255]^u[254]^u[239]^u[238]^u[223]^u[222]^u[207]^u[206]^u[191]^u[190]^u[175]^u[174]^u[159]^u[158]^u[143]^u[142]^u[127]^u[126]^u[111]^u[110]^u[95]^u[94]^u[79]^u[78]^u[63]^u[62]^u[47]^u[46]^u[31]^u[30]^u[15]^u[14],u[255]^u[254]^u[247]^u[246],u[255]^u[254]^u[247]^u[246]^u[127]^u[126]^u[119]^u[118],u[255]^u[254]^u[247]^u[246]^u[191]^u[190]^u[183]^u[182],u[255]^u[254]^u[247]^u[246]^u[191]^u[190]^u[183]^u[182]^u[127]^u[126]^u[119]^u[118]^u[63]^u[62]^u[55]^u[54],u[255]^u[254]^u[247]^u[246]^u[223]^u[222]^u[215]^u[214],u[255]^u[254]^u[247]^u[246]^u[223]^u[222]^u[215]^u[214]^u[127]^u[126]^u[119]^u[118]^u[95]^u[94]^u[87]^u[86],u[255]^u[254]^u[247]^u[246]^u[223]^u[222]^u[215]^u[214]^u[191]^u[190]^u[183]^u[182]^u[159]^u[158]^u[151]^u[150],u[255]^u[254]^u[247]^u[246]^u[223]^u[222]^u[215]^u[214]^u[191]^u[190]^u[183]^u[182]^u[159]^u[158]^u[151]^u[150]^u[127]^u[126]^u[119]^u[118]^u[95]^u[94]^u[87]^u[86]^u[63]^u[62]^u[55]^u[54]^u[31]^u[30]^u[23]^u[22],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[127]^u[126]^u[119]^u[118]^u[111]^u[110]^u[103]^u[102],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[191]^u[190]^u[183]^u[182]^u[175]^u[174]^u[167]^u[166],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[191]^u[190]^u[183]^u[182]^u[175]^u[174]^u[167]^u[166]^u[127]^u[126]^u[119]^u[118]^u[111]^u[110]^u[103]^u[102]^u[63]^u[62]^u[55]^u[54]^u[47]^u[46]^u[39]^u[38],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[223]^u[222]^u[215]^u[214]^u[207]^u[206]^u[199]^u[198],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[223]^u[222]^u[215]^u[214]^u[207]^u[206]^u[199]^u[198]^u[127]^u[126]^u[119]^u[118]^u[111]^u[110]^u[103]^u[102]^u[95]^u[94]^u[87]^u[86]^u[79]^u[78]^u[71]^u[70],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[223]^u[222]^u[215]^u[214]^u[207]^u[206]^u[199]^u[198]^u[191]^u[190]^u[183]^u[182]^u[175]^u[174]^u[167]^u[166]^u[159]^u[158]^u[151]^u[150]^u[143]^u[142]^u[135]^u[134],u[255]^u[254]^u[247]^u[246]^u[239]^u[238]^u[231]^u[230]^u[223]^u[222]^u[215]^u[214]^u[207]^u[206]^u[199]^u[198]^u[191]^u[190]^u[183]^u[182]^u[175]^u[174]^u[167]^u[166]^u[159]^u[158]^u[151]^u[150]^u[143]^u[142]^u[135]^u[134]^u[127]^u[126]^u[119]^u[118]^u[111]^u[110]^u[103]^u[102]^u[95]^u[94]^u[87]^u[86]^u[79]^u[78]^u[71]^u[70]^u[63]^u[62]^u[55]^u[54]^u[47]^u[46]^u[39]^u[38]^u[31]^u[30]^u[23]^u[22]^u[15]^u[14]^u[7]^u[6],u[255]^u[254]^u[251]^u[250],u[255]^u[254]^u[251]^u[250]^u[127]^u[126]^u[123]^u[122],u[255]^u[254]^u[251]^u[250]^u[191]^u[190]^u[187]^u[186],u[255]^u[254]^u[251]^u[250]^u[191]^u[190]^u[187]^u[186]^u[127]^u[126]^u[123]^u[122]^u[63]^u[62]^u[59]^u[58],u[255]^u[254]^u[251]^u[250]^u[223]^u[222]^u[219]^u[218],u[255]^u[254]^u[251]^u[250]^u[223]^u[222]^u[219]^u[218]^u[127]^u[126]^u[123]^u[122]^u[95]^u[94]^u[91]^u[90],u[255]^u[254]^u[251]^u[250]^u[223]^u[222]^u[219]^u[218]^u[191]^u[190]^u[187]^u[186]^u[159]^u[158]^u[155]^u[154],u[255]^u[254]^u[251]^u[250]^u[223]^u[222]^u[219]^u[218]^u[191]^u[190]^u[187]^u[186]^u[159]^u[158]^u[155]^u[154]^u[127]^u[126]^u[123]^u[122]^u[95]^u[94]^u[91]^u[90]^u[63]^u[62]^u[59]^u[58]^u[31]^u[30]^u[27]^u[26],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[127]^u[126]^u[123]^u[122]^u[111]^u[110]^u[107]^u[106],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[191]^u[190]^u[187]^u[186]^u[175]^u[174]^u[171]^u[170],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[191]^u[190]^u[187]^u[186]^u[175]^u[174]^u[171]^u[170]^u[127]^u[126]^u[123]^u[122]^u[111]^u[110]^u[107]^u[106]^u[63]^u[62]^u[59]^u[58]^u[47]^u[46]^u[43]^u[42],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[223]^u[222]^u[219]^u[218]^u[207]^u[206]^u[203]^u[202],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[223]^u[222]^u[219]^u[218]^u[207]^u[206]^u[203]^u[202]^u[127]^u[126]^u[123]^u[122]^u[111]^u[110]^u[107]^u[106]^u[95]^u[94]^u[91]^u[90]^u[79]^u[78]^u[75]^u[74],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[223]^u[222]^u[219]^u[218]^u[207]^u[206]^u[203]^u[202]^u[191]^u[190]^u[187]^u[186]^u[175]^u[174]^u[171]^u[170]^u[159]^u[158]^u[155]^u[154]^u[143]^u[142]^u[139]^u[138],u[255]^u[254]^u[251]^u[250]^u[239]^u[238]^u[235]^u[234]^u[223]^u[222]^u[219]^u[218]^u[207]^u[206]^u[203]^u[202]^u[191]^u[190]^u[187]^u[186]^u[175]^u[174]^u[171]^u[170]^u[159]^u[158]^u[155]^u[154]^u[143]^u[142]^u[139]^u[138]^u[127]^u[126]^u[123]^u[122]^u[111]^u[110]^u[107]^u[106]^u[95]^u[94]^u[91]^u[90]^u[79]^u[78]^u[75]^u[74]^u[63]^u[62]^u[59]^u[58]^u[47]^u[46]^u[43]^u[42]^u[31]^u[30]^u[27]^u[26]^u[15]^u[14]^u[11]^u[10],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[63]^u[62]^u[59]^u[58]^u[55]^u[54]^u[51]^u[50],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[95]^u[94]^u[91]^u[90]^u[87]^u[86]^u[83]^u[82],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[159]^u[158]^u[155]^u[154]^u[151]^u[150]^u[147]^u[146],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[159]^u[158]^u[155]^u[154]^u[151]^u[150]^u[147]^u[146]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[95]^u[94]^u[91]^u[90]^u[87]^u[86]^u[83]^u[82]^u[63]^u[62]^u[59]^u[58]^u[55]^u[54]^u[51]^u[50]^u[31]^u[30]^u[27]^u[26]^u[23]^u[22]^u[19]^u[18],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[111]^u[110]^u[107]^u[106]^u[103]^u[102]^u[99]^u[98],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[175]^u[174]^u[171]^u[170]^u[167]^u[166]^u[163]^u[162],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[175]^u[174]^u[171]^u[170]^u[167]^u[166]^u[163]^u[162]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[111]^u[110]^u[107]^u[106]^u[103]^u[102]^u[99]^u[98]^u[63]^u[62]^u[59]^u[58]^u[55]^u[54]^u[51]^u[50]^u[47]^u[46]^u[43]^u[42]^u[39]^u[38]^u[35]^u[34],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[207]^u[206]^u[203]^u[202]^u[199]^u[198]^u[195]^u[194],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[207]^u[206]^u[203]^u[202]^u[199]^u[198]^u[195]^u[194]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[111]^u[110]^u[107]^u[106]^u[103]^u[102]^u[99]^u[98]^u[95]^u[94]^u[91]^u[90]^u[87]^u[86]^u[83]^u[82]^u[79]^u[78]^u[75]^u[74]^u[71]^u[70]^u[67]^u[66],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[207]^u[206]^u[203]^u[202]^u[199]^u[198]^u[195]^u[194]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[175]^u[174]^u[171]^u[170]^u[167]^u[166]^u[163]^u[162]^u[159]^u[158]^u[155]^u[154]^u[151]^u[150]^u[147]^u[146]^u[143]^u[142]^u[139]^u[138]^u[135]^u[134]^u[131]^u[130],u[255]^u[254]^u[251]^u[250]^u[247]^u[246]^u[243]^u[242]^u[239]^u[238]^u[235]^u[234]^u[231]^u[230]^u[227]^u[226]^u[223]^u[222]^u[219]^u[218]^u[215]^u[214]^u[211]^u[210]^u[207]^u[206]^u[203]^u[202]^u[199]^u[198]^u[195]^u[194]^u[191]^u[190]^u[187]^u[186]^u[183]^u[182]^u[179]^u[178]^u[175]^u[174]^u[171]^u[170]^u[167]^u[166]^u[163]^u[162]^u[159]^u[158]^u[155]^u[154]^u[151]^u[150]^u[147]^u[146]^u[143]^u[142]^u[139]^u[138]^u[135]^u[134]^u[131]^u[130]^u[127]^u[126]^u[123]^u[122]^u[119]^u[118]^u[115]^u[114]^u[111]^u[110]^u[107]^u[106]^u[103]^u[102]^u[99]^u[98]^u[95]^u[94]^u[91]^u[90]^u[87]^u[86]^u[83]^u[82]^u[79]^u[78]^u[75]^u[74]^u[71]^u[70]^u[67]^u[66]^u[63]^u[62]^u[59]^u[58]^u[55]^u[54]^u[51]^u[50]^u[47]^u[46]^u[43]^u[42]^u[39]^u[38]^u[35]^u[34]^u[31]^u[30]^u[27]^u[26]^u[23]^u[22]^u[19]^u[18]^u[15]^u[14]^u[11]^u[10]^u[7]^u[6]^u[3]^u[2],u[255]^u[254]^u[253]^u[252],u[255]^u[254]^u[253]^u[252]^u[127]^u[126]^u[125]^u[124],u[255]^u[254]^u[253]^u[252]^u[191]^u[190]^u[189]^u[188],u[255]^u[254]^u[253]^u[252]^u[191]^u[190]^u[189]^u[188]^u[127]^u[126]^u[125]^u[124]^u[63]^u[62]^u[61]^u[60],u[255]^u[254]^u[253]^u[252]^u[223]^u[222]^u[221]^u[220],u[255]^u[254]^u[253]^u[252]^u[223]^u[222]^u[221]^u[220]^u[127]^u[126]^u[125]^u[124]^u[95]^u[94]^u[93]^u[92],u[255]^u[254]^u[253]^u[252]^u[223]^u[222]^u[221]^u[220]^u[191]^u[190]^u[189]^u[188]^u[159]^u[158]^u[157]^u[156],u[255]^u[254]^u[253]^u[252]^u[223]^u[222]^u[221]^u[220]^u[191]^u[190]^u[189]^u[188]^u[159]^u[158]^u[157]^u[156]^u[127]^u[126]^u[125]^u[124]^u[95]^u[94]^u[93]^u[92]^u[63]^u[62]^u[61]^u[60]^u[31]^u[30]^u[29]^u[28],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[127]^u[126]^u[125]^u[124]^u[111]^u[110]^u[109]^u[108],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[191]^u[190]^u[189]^u[188]^u[175]^u[174]^u[173]^u[172],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[191]^u[190]^u[189]^u[188]^u[175]^u[174]^u[173]^u[172]^u[127]^u[126]^u[125]^u[124]^u[111]^u[110]^u[109]^u[108]^u[63]^u[62]^u[61]^u[60]^u[47]^u[46]^u[45]^u[44],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[223]^u[222]^u[221]^u[220]^u[207]^u[206]^u[205]^u[204],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[223]^u[222]^u[221]^u[220]^u[207]^u[206]^u[205]^u[204]^u[127]^u[126]^u[125]^u[124]^u[111]^u[110]^u[109]^u[108]^u[95]^u[94]^u[93]^u[92]^u[79]^u[78]^u[77]^u[76],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[223]^u[222]^u[221]^u[220]^u[207]^u[206]^u[205]^u[204]^u[191]^u[190]^u[189]^u[188]^u[175]^u[174]^u[173]^u[172]^u[159]^u[158]^u[157]^u[156]^u[143]^u[142]^u[141]^u[140],u[255]^u[254]^u[253]^u[252]^u[239]^u[238]^u[237]^u[236]^u[223]^u[222]^u[221]^u[220]^u[207]^u[206]^u[205]^u[204]^u[191]^u[190]^u[189]^u[188]^u[175]^u[174]^u[173]^u[172]^u[159]^u[158]^u[157]^u[156]^u[143]^u[142]^u[141]^u[140]^u[127]^u[126]^u[125]^u[124]^u[111]^u[110]^u[109]^u[108]^u[95]^u[94]^u[93]^u[92]^u[79]^u[78]^u[77]^u[76]^u[63]^u[62]^u[61]^u[60]^u[47]^u[46]^u[45]^u[44]^u[31]^u[30]^u[29]^u[28]^u[15]^u[14]^u[13]^u[12],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[63]^u[62]^u[61]^u[60]^u[55]^u[54]^u[53]^u[52],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[95]^u[94]^u[93]^u[92]^u[87]^u[86]^u[85]^u[84],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[159]^u[158]^u[157]^u[156]^u[151]^u[150]^u[149]^u[148],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[159]^u[158]^u[157]^u[156]^u[151]^u[150]^u[149]^u[148]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[95]^u[94]^u[93]^u[92]^u[87]^u[86]^u[85]^u[84]^u[63]^u[62]^u[61]^u[60]^u[55]^u[54]^u[53]^u[52]^u[31]^u[30]^u[29]^u[28]^u[23]^u[22]^u[21]^u[20],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[111]^u[110]^u[109]^u[108]^u[103]^u[102]^u[101]^u[100],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[175]^u[174]^u[173]^u[172]^u[167]^u[166]^u[165]^u[164],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[175]^u[174]^u[173]^u[172]^u[167]^u[166]^u[165]^u[164]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[111]^u[110]^u[109]^u[108]^u[103]^u[102]^u[101]^u[100]^u[63]^u[62]^u[61]^u[60]^u[55]^u[54]^u[53]^u[52]^u[47]^u[46]^u[45]^u[44]^u[39]^u[38]^u[37]^u[36],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[207]^u[206]^u[205]^u[204]^u[199]^u[198]^u[197]^u[196],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[207]^u[206]^u[205]^u[204]^u[199]^u[198]^u[197]^u[196]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[111]^u[110]^u[109]^u[108]^u[103]^u[102]^u[101]^u[100]^u[95]^u[94]^u[93]^u[92]^u[87]^u[86]^u[85]^u[84]^u[79]^u[78]^u[77]^u[76]^u[71]^u[70]^u[69]^u[68],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[207]^u[206]^u[205]^u[204]^u[199]^u[198]^u[197]^u[196]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[175]^u[174]^u[173]^u[172]^u[167]^u[166]^u[165]^u[164]^u[159]^u[158]^u[157]^u[156]^u[151]^u[150]^u[149]^u[148]^u[143]^u[142]^u[141]^u[140]^u[135]^u[134]^u[133]^u[132],u[255]^u[254]^u[253]^u[252]^u[247]^u[246]^u[245]^u[244]^u[239]^u[238]^u[237]^u[236]^u[231]^u[230]^u[229]^u[228]^u[223]^u[222]^u[221]^u[220]^u[215]^u[214]^u[213]^u[212]^u[207]^u[206]^u[205]^u[204]^u[199]^u[198]^u[197]^u[196]^u[191]^u[190]^u[189]^u[188]^u[183]^u[182]^u[181]^u[180]^u[175]^u[174]^u[173]^u[172]^u[167]^u[166]^u[165]^u[164]^u[159]^u[158]^u[157]^u[156]^u[151]^u[150]^u[149]^u[148]^u[143]^u[142]^u[141]^u[140]^u[135]^u[134]^u[133]^u[132]^u[127]^u[126]^u[125]^u[124]^u[119]^u[118]^u[117]^u[116]^u[111]^u[110]^u[109]^u[108]^u[103]^u[102]^u[101]^u[100]^u[95]^u[94]^u[93]^u[92]^u[87]^u[86]^u[85]^u[84]^u[79]^u[78]^u[77]^u[76]^u[71]^u[70]^u[69]^u[68]^u[63]^u[62]^u[61]^u[60]^u[55]^u[54]^u[53]^u[52]^u[47]^u[46]^u[45]^u[44]^u[39]^u[38]^u[37]^u[36]^u[31]^u[30]^u[29]^u[28]^u[23]^u[22]^u[21]^u[20]^u[15]^u[14]^u[13]^u[12]^u[7]^u[6]^u[5]^u[4],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[79]^u[78]^u[77]^u[76]^u[75]^u[74]^u[73]^u[72],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[143]^u[142]^u[141]^u[140]^u[139]^u[138]^u[137]^u[136],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[143]^u[142]^u[141]^u[140]^u[139]^u[138]^u[137]^u[136]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[79]^u[78]^u[77]^u[76]^u[75]^u[74]^u[73]^u[72]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[87]^u[86]^u[85]^u[84]^u[83]^u[82]^u[81]^u[80],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[151]^u[150]^u[149]^u[148]^u[147]^u[146]^u[145]^u[144],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[151]^u[150]^u[149]^u[148]^u[147]^u[146]^u[145]^u[144]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[87]^u[86]^u[85]^u[84]^u[83]^u[82]^u[81]^u[80]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[103]^u[102]^u[101]^u[100]^u[99]^u[98]^u[97]^u[96],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[167]^u[166]^u[165]^u[164]^u[163]^u[162]^u[161]^u[160],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[167]^u[166]^u[165]^u[164]^u[163]^u[162]^u[161]^u[160]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[103]^u[102]^u[101]^u[100]^u[99]^u[98]^u[97]^u[96]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[199]^u[198]^u[197]^u[196]^u[195]^u[194]^u[193]^u[192],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[199]^u[198]^u[197]^u[196]^u[195]^u[194]^u[193]^u[192]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[103]^u[102]^u[101]^u[100]^u[99]^u[98]^u[97]^u[96]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[87]^u[86]^u[85]^u[84]^u[83]^u[82]^u[81]^u[80]^u[79]^u[78]^u[77]^u[76]^u[75]^u[74]^u[73]^u[72]^u[71]^u[70]^u[69]^u[68]^u[67]^u[66]^u[65]^u[64],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[199]^u[198]^u[197]^u[196]^u[195]^u[194]^u[193]^u[192]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[167]^u[166]^u[165]^u[164]^u[163]^u[162]^u[161]^u[160]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[151]^u[150]^u[149]^u[148]^u[147]^u[146]^u[145]^u[144]^u[143]^u[142]^u[141]^u[140]^u[139]^u[138]^u[137]^u[136]^u[135]^u[134]^u[133]^u[132]^u[131]^u[130]^u[129]^u[128],u[255]^u[254]^u[253]^u[252]^u[251]^u[250]^u[249]^u[248]^u[247]^u[246]^u[245]^u[244]^u[243]^u[242]^u[241]^u[240]^u[239]^u[238]^u[237]^u[236]^u[235]^u[234]^u[233]^u[232]^u[231]^u[230]^u[229]^u[228]^u[227]^u[226]^u[225]^u[224]^u[223]^u[222]^u[221]^u[220]^u[219]^u[218]^u[217]^u[216]^u[215]^u[214]^u[213]^u[212]^u[211]^u[210]^u[209]^u[208]^u[207]^u[206]^u[205]^u[204]^u[203]^u[202]^u[201]^u[200]^u[199]^u[198]^u[197]^u[196]^u[195]^u[194]^u[193]^u[192]^u[191]^u[190]^u[189]^u[188]^u[187]^u[186]^u[185]^u[184]^u[183]^u[182]^u[181]^u[180]^u[179]^u[178]^u[177]^u[176]^u[175]^u[174]^u[173]^u[172]^u[171]^u[170]^u[169]^u[168]^u[167]^u[166]^u[165]^u[164]^u[163]^u[162]^u[161]^u[160]^u[159]^u[158]^u[157]^u[156]^u[155]^u[154]^u[153]^u[152]^u[151]^u[150]^u[149]^u[148]^u[147]^u[146]^u[145]^u[144]^u[143]^u[142]^u[141]^u[140]^u[139]^u[138]^u[137]^u[136]^u[135]^u[134]^u[133]^u[132]^u[131]^u[130]^u[129]^u[128]^u[127]^u[126]^u[125]^u[124]^u[123]^u[122]^u[121]^u[120]^u[119]^u[118]^u[117]^u[116]^u[115]^u[114]^u[113]^u[112]^u[111]^u[110]^u[109]^u[108]^u[107]^u[106]^u[105]^u[104]^u[103]^u[102]^u[101]^u[100]^u[99]^u[98]^u[97]^u[96]^u[95]^u[94]^u[93]^u[92]^u[91]^u[90]^u[89]^u[88]^u[87]^u[86]^u[85]^u[84]^u[83]^u[82]^u[81]^u[80]^u[79]^u[78]^u[77]^u[76]^u[75]^u[74]^u[73]^u[72]^u[71]^u[70]^u[69]^u[68]^u[67]^u[66]^u[65]^u[64]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0]};
assign usum_128 = {usum_256[255],usum_256[253],usum_256[251],usum_256[249],usum_256[247],usum_256[245],usum_256[243],usum_256[241],usum_256[239],usum_256[237],usum_256[235],usum_256[233],usum_256[231],usum_256[229],usum_256[227],usum_256[225],usum_256[223],usum_256[221],usum_256[219],usum_256[217],usum_256[215],usum_256[213],usum_256[211],usum_256[209],usum_256[207],usum_256[205],usum_256[203],usum_256[201],usum_256[199],usum_256[197],usum_256[195],usum_256[193],usum_256[191],usum_256[189],usum_256[187],usum_256[185],usum_256[183],usum_256[181],usum_256[179],usum_256[177],usum_256[175],usum_256[173],usum_256[171],usum_256[169],usum_256[167],usum_256[165],usum_256[163],usum_256[161],usum_256[159],usum_256[157],usum_256[155],usum_256[153],usum_256[151],usum_256[149],usum_256[147],usum_256[145],usum_256[143],usum_256[141],usum_256[139],usum_256[137],usum_256[135],usum_256[133],usum_256[131],usum_256[129],usum_256[127],usum_256[125],usum_256[123],usum_256[121],usum_256[119],usum_256[117],usum_256[115],usum_256[113],usum_256[111],usum_256[109],usum_256[107],usum_256[105],usum_256[103],usum_256[101],usum_256[99],usum_256[97],usum_256[95],usum_256[93],usum_256[91],usum_256[89],usum_256[87],usum_256[85],usum_256[83],usum_256[81],usum_256[79],usum_256[77],usum_256[75],usum_256[73],usum_256[71],usum_256[69],usum_256[67],usum_256[65],usum_256[63],usum_256[61],usum_256[59],usum_256[57],usum_256[55],usum_256[53],usum_256[51],usum_256[49],usum_256[47],usum_256[45],usum_256[43],usum_256[41],usum_256[39],usum_256[37],usum_256[35],usum_256[33],usum_256[31],usum_256[29],usum_256[27],usum_256[25],usum_256[23],usum_256[21],usum_256[19],usum_256[17],usum_256[15],usum_256[13],usum_256[11],usum_256[9],usum_256[7],usum_256[5],usum_256[3],usum_256[1]};
assign usum_64  = {usum_256[255],usum_256[251],usum_256[247],usum_256[243],usum_256[239],usum_256[235],usum_256[231],usum_256[227],usum_256[223],usum_256[219],usum_256[215],usum_256[211],usum_256[207],usum_256[203],usum_256[199],usum_256[195],usum_256[191],usum_256[187],usum_256[183],usum_256[179],usum_256[175],usum_256[171],usum_256[167],usum_256[163],usum_256[159],usum_256[155],usum_256[151],usum_256[147],usum_256[143],usum_256[139],usum_256[135],usum_256[131],usum_256[127],usum_256[123],usum_256[119],usum_256[115],usum_256[111],usum_256[107],usum_256[103],usum_256[99],usum_256[95],usum_256[91],usum_256[87],usum_256[83],usum_256[79],usum_256[75],usum_256[71],usum_256[67],usum_256[63],usum_256[59],usum_256[55],usum_256[51],usum_256[47],usum_256[43],usum_256[39],usum_256[35],usum_256[31],usum_256[27],usum_256[23],usum_256[19],usum_256[15],usum_256[11],usum_256[7],usum_256[3]};
assign usum_32  = {usum_256[255],usum_256[247],usum_256[239],usum_256[231],usum_256[223],usum_256[215],usum_256[207],usum_256[199],usum_256[191],usum_256[183],usum_256[175],usum_256[167],usum_256[159],usum_256[151],usum_256[143],usum_256[135],usum_256[127],usum_256[119],usum_256[111],usum_256[103],usum_256[95],usum_256[87],usum_256[79],usum_256[71],usum_256[63],usum_256[55],usum_256[47],usum_256[39],usum_256[31],usum_256[23],usum_256[15],usum_256[7]};
assign usum_16  = {usum_256[255],usum_256[239],usum_256[223],usum_256[207],usum_256[191],usum_256[175],usum_256[159],usum_256[143],usum_256[127],usum_256[111],usum_256[95],usum_256[79],usum_256[63],usum_256[47],usum_256[31],usum_256[15]};
assign usum_8   = {usum_256[255],usum_256[223],usum_256[191],usum_256[159],usum_256[127],usum_256[95],usum_256[63],usum_256[31]};
assign usum_4   = {usum_256[255],usum_256[191],usum_256[127],usum_256[63]};
assign usum_2   = {usum_256[255],usum_256[127]};

always @(posedge clk or negedge rst_n) begin
	if(!rst_n)
		u <= 0;
	else if(state==DONE)
		u <= 0;
	else if(state==DECODE && counter[0]==0 && counter<N)
		u <= {pnode_N,u[255:2]};
	else
		u <= u;
end

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		usum2   <= 0;
		usum4   <= 0;
		usum8   <= 0;
		usum16  <= 0;
		usum32  <= 0;
		usum64  <= 0;
		usum128 <= 0;
		usum256 <= 0;
	end else if(state==DONE) begin
		usum2   <= 0;
		usum4   <= 0;
		usum8   <= 0;
		usum16  <= 0;
		usum32  <= 0;
		usum64  <= 0;
		usum128 <= 0;
		usum256 <= 0;
	end else if(state==DECODE && counter[0]==1 && counter<N-2) begin
		usum2   <= (~usum_counter_minus[0] && usum_counter[0]) ? usum_2   : usum2;
		usum4   <= (~usum_counter_minus[1] && usum_counter[1]) ? usum_4   : usum4;
		usum8   <= (~usum_counter_minus[2] && usum_counter[2]) ? usum_8   : usum8;
		usum16  <= (~usum_counter_minus[3] && usum_counter[3]) ? usum_16  : usum16;
		usum32  <= (~usum_counter_minus[4] && usum_counter[4]) ? usum_32  : usum32;
		usum64  <= (~usum_counter_minus[5] && usum_counter[5]) ? usum_64  : usum64;
		usum128 <= (~usum_counter_minus[6] && usum_counter[6]) ? usum_128 : usum128;
		usum256 <= (~usum_counter_minus[7] && usum_counter[7]) ? usum_256 : usum256;
	end else begin
		usum2   <= usum2;
		usum4   <= usum4;
		usum8   <= usum8;
		usum16  <= usum16;
		usum32  <= usum32;
		usum64  <= usum64;
		usum128 <= usum128;
		usum256 <= usum256;
	end
end

assign input1_128 = PE(PE(PE(PE(PE(PE(LLR[1],LLR[65],u_counter[5],usum64[0]),PE(LLR[33],LLR[97],u_counter[5],usum64[1]),u_counter[4],usum32[0]),PE(PE(LLR[17],LLR[81],u_counter[5],usum64[2]),PE(LLR[49],LLR[113],u_counter[5],usum64[3]),u_counter[4],usum32[1]),u_counter[3],usum16[0]),PE(PE(PE(LLR[9],LLR[73],u_counter[5],usum64[4]),PE(LLR[41],LLR[105],u_counter[5],usum64[5]),u_counter[4],usum32[2]),PE(PE(LLR[25],LLR[89],u_counter[5],usum64[6]),PE(LLR[57],LLR[121],u_counter[5],usum64[7]),u_counter[4],usum32[3]),u_counter[3],usum16[1]),u_counter[2],usum8[0]),PE(PE(PE(PE(LLR[5],LLR[69],u_counter[5],usum64[8]),PE(LLR[37],LLR[101],u_counter[5],usum64[9]),u_counter[4],usum32[4]),PE(PE(LLR[21],LLR[85],u_counter[5],usum64[10]),PE(LLR[53],LLR[117],u_counter[5],usum64[11]),u_counter[4],usum32[5]),u_counter[3],usum16[2]),PE(PE(PE(LLR[13],LLR[77],u_counter[5],usum64[12]),PE(LLR[45],LLR[109],u_counter[5],usum64[13]),u_counter[4],usum32[6]),PE(PE(LLR[29],LLR[93],u_counter[5],usum64[14]),PE(LLR[61],LLR[125],u_counter[5],usum64[15]),u_counter[4],usum32[7]),u_counter[3],usum16[3]),u_counter[2],usum8[1]),u_counter[1],usum4[0]),PE(PE(PE(PE(PE(LLR[3],LLR[67],u_counter[5],usum64[16]),PE(LLR[35],LLR[99],u_counter[5],usum64[17]),u_counter[4],usum32[8]),PE(PE(LLR[19],LLR[83],u_counter[5],usum64[18]),PE(LLR[51],LLR[115],u_counter[5],usum64[19]),u_counter[4],usum32[9]),u_counter[3],usum16[4]),PE(PE(PE(LLR[11],LLR[75],u_counter[5],usum64[20]),PE(LLR[43],LLR[107],u_counter[5],usum64[21]),u_counter[4],usum32[10]),PE(PE(LLR[27],LLR[91],u_counter[5],usum64[22]),PE(LLR[59],LLR[123],u_counter[5],usum64[23]),u_counter[4],usum32[11]),u_counter[3],usum16[5]),u_counter[2],usum8[2]),PE(PE(PE(PE(LLR[7],LLR[71],u_counter[5],usum64[24]),PE(LLR[39],LLR[103],u_counter[5],usum64[25]),u_counter[4],usum32[12]),PE(PE(LLR[23],LLR[87],u_counter[5],usum64[26]),PE(LLR[55],LLR[119],u_counter[5],usum64[27]),u_counter[4],usum32[13]),u_counter[3],usum16[6]),PE(PE(PE(LLR[15],LLR[79],u_counter[5],usum64[28]),PE(LLR[47],LLR[111],u_counter[5],usum64[29]),u_counter[4],usum32[14]),PE(PE(LLR[31],LLR[95],u_counter[5],usum64[30]),PE(LLR[63],LLR[127],u_counter[5],usum64[31]),u_counter[4],usum32[15]),u_counter[3],usum16[7]),u_counter[2],usum8[3]),u_counter[1],usum4[1]),u_counter[0],usum2[0]);
assign input2_128 = PE(PE(PE(PE(PE(PE(LLR[2],LLR[66],u_counter[5],usum64[32]),PE(LLR[34],LLR[98],u_counter[5],usum64[33]),u_counter[4],usum32[16]),PE(PE(LLR[18],LLR[82],u_counter[5],usum64[34]),PE(LLR[50],LLR[114],u_counter[5],usum64[35]),u_counter[4],usum32[17]),u_counter[3],usum16[8]),PE(PE(PE(LLR[10],LLR[74],u_counter[5],usum64[36]),PE(LLR[42],LLR[106],u_counter[5],usum64[37]),u_counter[4],usum32[18]),PE(PE(LLR[26],LLR[90],u_counter[5],usum64[38]),PE(LLR[58],LLR[122],u_counter[5],usum64[39]),u_counter[4],usum32[19]),u_counter[3],usum16[9]),u_counter[2],usum8[4]),PE(PE(PE(PE(LLR[6],LLR[70],u_counter[5],usum64[40]),PE(LLR[38],LLR[102],u_counter[5],usum64[41]),u_counter[4],usum32[20]),PE(PE(LLR[22],LLR[86],u_counter[5],usum64[42]),PE(LLR[54],LLR[118],u_counter[5],usum64[43]),u_counter[4],usum32[21]),u_counter[3],usum16[10]),PE(PE(PE(LLR[14],LLR[78],u_counter[5],usum64[44]),PE(LLR[46],LLR[110],u_counter[5],usum64[45]),u_counter[4],usum32[22]),PE(PE(LLR[30],LLR[94],u_counter[5],usum64[46]),PE(LLR[62],LLR[126],u_counter[5],usum64[47]),u_counter[4],usum32[23]),u_counter[3],usum16[11]),u_counter[2],usum8[5]),u_counter[1],usum4[2]),PE(PE(PE(PE(PE(LLR[4],LLR[68],u_counter[5],usum64[48]),PE(LLR[36],LLR[100],u_counter[5],usum64[49]),u_counter[4],usum32[24]),PE(PE(LLR[20],LLR[84],u_counter[5],usum64[50]),PE(LLR[52],LLR[116],u_counter[5],usum64[51]),u_counter[4],usum32[25]),u_counter[3],usum16[12]),PE(PE(PE(LLR[12],LLR[76],u_counter[5],usum64[52]),PE(LLR[44],LLR[108],u_counter[5],usum64[53]),u_counter[4],usum32[26]),PE(PE(LLR[28],LLR[92],u_counter[5],usum64[54]),PE(LLR[60],LLR[124],u_counter[5],usum64[55]),u_counter[4],usum32[27]),u_counter[3],usum16[13]),u_counter[2],usum8[6]),PE(PE(PE(PE(LLR[8],LLR[72],u_counter[5],usum64[56]),PE(LLR[40],LLR[104],u_counter[5],usum64[57]),u_counter[4],usum32[28]),PE(PE(LLR[24],LLR[88],u_counter[5],usum64[58]),PE(LLR[56],LLR[120],u_counter[5],usum64[59]),u_counter[4],usum32[29]),u_counter[3],usum16[14]),PE(PE(PE(LLR[16],LLR[80],u_counter[5],usum64[60]),PE(LLR[48],LLR[112],u_counter[5],usum64[61]),u_counter[4],usum32[30]),PE(PE(LLR[32],LLR[96],u_counter[5],usum64[62]),PE(LLR[64],LLR[128],u_counter[5],usum64[63]),u_counter[4],usum32[31]),u_counter[3],usum16[15]),u_counter[2],usum8[7]),u_counter[1],usum4[3]),u_counter[0],usum2[1]);
assign input1_256 = PE(PE(PE(PE(PE(PE(PE(LLR[1],LLR[129],u_counter[6],usum128[0]),PE(LLR[65],LLR[193],u_counter[6],usum128[1]),u_counter[5],usum64[0]),PE(PE(LLR[33],LLR[161],u_counter[6],usum128[2]),PE(LLR[97],LLR[225],u_counter[6],usum128[3]),u_counter[5],usum64[1]),u_counter[4],usum32[0]),PE(PE(PE(LLR[17],LLR[145],u_counter[6],usum128[4]),PE(LLR[81],LLR[209],u_counter[6],usum128[5]),u_counter[5],usum64[2]),PE(PE(LLR[49],LLR[177],u_counter[6],usum128[6]),PE(LLR[113],LLR[241],u_counter[6],usum128[7]),u_counter[5],usum64[3]),u_counter[4],usum32[1]),u_counter[3],usum16[0]),PE(PE(PE(PE(LLR[9],LLR[137],u_counter[6],usum128[8]),PE(LLR[73],LLR[201],u_counter[6],usum128[9]),u_counter[5],usum64[4]),PE(PE(LLR[41],LLR[169],u_counter[6],usum128[10]),PE(LLR[105],LLR[233],u_counter[6],usum128[11]),u_counter[5],usum64[5]),u_counter[4],usum32[2]),PE(PE(PE(LLR[25],LLR[153],u_counter[6],usum128[12]),PE(LLR[89],LLR[217],u_counter[6],usum128[13]),u_counter[5],usum64[6]),PE(PE(LLR[57],LLR[185],u_counter[6],usum128[14]),PE(LLR[121],LLR[249],u_counter[6],usum128[15]),u_counter[5],usum64[7]),u_counter[4],usum32[3]),u_counter[3],usum16[1]),u_counter[2],usum8[0]),PE(PE(PE(PE(PE(LLR[5],LLR[133],u_counter[6],usum128[16]),PE(LLR[69],LLR[197],u_counter[6],usum128[17]),u_counter[5],usum64[8]),PE(PE(LLR[37],LLR[165],u_counter[6],usum128[18]),PE(LLR[101],LLR[229],u_counter[6],usum128[19]),u_counter[5],usum64[9]),u_counter[4],usum32[4]),PE(PE(PE(LLR[21],LLR[149],u_counter[6],usum128[20]),PE(LLR[85],LLR[213],u_counter[6],usum128[21]),u_counter[5],usum64[10]),PE(PE(LLR[53],LLR[181],u_counter[6],usum128[22]),PE(LLR[117],LLR[245],u_counter[6],usum128[23]),u_counter[5],usum64[11]),u_counter[4],usum32[5]),u_counter[3],usum16[2]),PE(PE(PE(PE(LLR[13],LLR[141],u_counter[6],usum128[24]),PE(LLR[77],LLR[205],u_counter[6],usum128[25]),u_counter[5],usum64[12]),PE(PE(LLR[45],LLR[173],u_counter[6],usum128[26]),PE(LLR[109],LLR[237],u_counter[6],usum128[27]),u_counter[5],usum64[13]),u_counter[4],usum32[6]),PE(PE(PE(LLR[29],LLR[157],u_counter[6],usum128[28]),PE(LLR[93],LLR[221],u_counter[6],usum128[29]),u_counter[5],usum64[14]),PE(PE(LLR[61],LLR[189],u_counter[6],usum128[30]),PE(LLR[125],LLR[253],u_counter[6],usum128[31]),u_counter[5],usum64[15]),u_counter[4],usum32[7]),u_counter[3],usum16[3]),u_counter[2],usum8[1]),u_counter[1],usum4[0]),PE(PE(PE(PE(PE(PE(LLR[3],LLR[131],u_counter[6],usum128[32]),PE(LLR[67],LLR[195],u_counter[6],usum128[33]),u_counter[5],usum64[16]),PE(PE(LLR[35],LLR[163],u_counter[6],usum128[34]),PE(LLR[99],LLR[227],u_counter[6],usum128[35]),u_counter[5],usum64[17]),u_counter[4],usum32[8]),PE(PE(PE(LLR[19],LLR[147],u_counter[6],usum128[36]),PE(LLR[83],LLR[211],u_counter[6],usum128[37]),u_counter[5],usum64[18]),PE(PE(LLR[51],LLR[179],u_counter[6],usum128[38]),PE(LLR[115],LLR[243],u_counter[6],usum128[39]),u_counter[5],usum64[19]),u_counter[4],usum32[9]),u_counter[3],usum16[4]),PE(PE(PE(PE(LLR[11],LLR[139],u_counter[6],usum128[40]),PE(LLR[75],LLR[203],u_counter[6],usum128[41]),u_counter[5],usum64[20]),PE(PE(LLR[43],LLR[171],u_counter[6],usum128[42]),PE(LLR[107],LLR[235],u_counter[6],usum128[43]),u_counter[5],usum64[21]),u_counter[4],usum32[10]),PE(PE(PE(LLR[27],LLR[155],u_counter[6],usum128[44]),PE(LLR[91],LLR[219],u_counter[6],usum128[45]),u_counter[5],usum64[22]),PE(PE(LLR[59],LLR[187],u_counter[6],usum128[46]),PE(LLR[123],LLR[251],u_counter[6],usum128[47]),u_counter[5],usum64[23]),u_counter[4],usum32[11]),u_counter[3],usum16[5]),u_counter[2],usum8[2]),PE(PE(PE(PE(PE(LLR[7],LLR[135],u_counter[6],usum128[48]),PE(LLR[71],LLR[199],u_counter[6],usum128[49]),u_counter[5],usum64[24]),PE(PE(LLR[39],LLR[167],u_counter[6],usum128[50]),PE(LLR[103],LLR[231],u_counter[6],usum128[51]),u_counter[5],usum64[25]),u_counter[4],usum32[12]),PE(PE(PE(LLR[23],LLR[151],u_counter[6],usum128[52]),PE(LLR[87],LLR[215],u_counter[6],usum128[53]),u_counter[5],usum64[26]),PE(PE(LLR[55],LLR[183],u_counter[6],usum128[54]),PE(LLR[119],LLR[247],u_counter[6],usum128[55]),u_counter[5],usum64[27]),u_counter[4],usum32[13]),u_counter[3],usum16[6]),PE(PE(PE(PE(LLR[15],LLR[143],u_counter[6],usum128[56]),PE(LLR[79],LLR[207],u_counter[6],usum128[57]),u_counter[5],usum64[28]),PE(PE(LLR[47],LLR[175],u_counter[6],usum128[58]),PE(LLR[111],LLR[239],u_counter[6],usum128[59]),u_counter[5],usum64[29]),u_counter[4],usum32[14]),PE(PE(PE(LLR[31],LLR[159],u_counter[6],usum128[60]),PE(LLR[95],LLR[223],u_counter[6],usum128[61]),u_counter[5],usum64[30]),PE(PE(LLR[63],LLR[191],u_counter[6],usum128[62]),PE(LLR[127],LLR[255],u_counter[6],usum128[63]),u_counter[5],usum64[31]),u_counter[4],usum32[15]),u_counter[3],usum16[7]),u_counter[2],usum8[3]),u_counter[1],usum4[1]),u_counter[0],usum2[0]);
assign input2_256 = PE(PE(PE(PE(PE(PE(PE(LLR[2],LLR[130],u_counter[6],usum128[64]),PE(LLR[66],LLR[194],u_counter[6],usum128[65]),u_counter[5],usum64[32]),PE(PE(LLR[34],LLR[162],u_counter[6],usum128[66]),PE(LLR[98],LLR[226],u_counter[6],usum128[67]),u_counter[5],usum64[33]),u_counter[4],usum32[16]),PE(PE(PE(LLR[18],LLR[146],u_counter[6],usum128[68]),PE(LLR[82],LLR[210],u_counter[6],usum128[69]),u_counter[5],usum64[34]),PE(PE(LLR[50],LLR[178],u_counter[6],usum128[70]),PE(LLR[114],LLR[242],u_counter[6],usum128[71]),u_counter[5],usum64[35]),u_counter[4],usum32[17]),u_counter[3],usum16[8]),PE(PE(PE(PE(LLR[10],LLR[138],u_counter[6],usum128[72]),PE(LLR[74],LLR[202],u_counter[6],usum128[73]),u_counter[5],usum64[36]),PE(PE(LLR[42],LLR[170],u_counter[6],usum128[74]),PE(LLR[106],LLR[234],u_counter[6],usum128[75]),u_counter[5],usum64[37]),u_counter[4],usum32[18]),PE(PE(PE(LLR[26],LLR[154],u_counter[6],usum128[76]),PE(LLR[90],LLR[218],u_counter[6],usum128[77]),u_counter[5],usum64[38]),PE(PE(LLR[58],LLR[186],u_counter[6],usum128[78]),PE(LLR[122],LLR[250],u_counter[6],usum128[79]),u_counter[5],usum64[39]),u_counter[4],usum32[19]),u_counter[3],usum16[9]),u_counter[2],usum8[4]),PE(PE(PE(PE(PE(LLR[6],LLR[134],u_counter[6],usum128[80]),PE(LLR[70],LLR[198],u_counter[6],usum128[81]),u_counter[5],usum64[40]),PE(PE(LLR[38],LLR[166],u_counter[6],usum128[82]),PE(LLR[102],LLR[230],u_counter[6],usum128[83]),u_counter[5],usum64[41]),u_counter[4],usum32[20]),PE(PE(PE(LLR[22],LLR[150],u_counter[6],usum128[84]),PE(LLR[86],LLR[214],u_counter[6],usum128[85]),u_counter[5],usum64[42]),PE(PE(LLR[54],LLR[182],u_counter[6],usum128[86]),PE(LLR[118],LLR[246],u_counter[6],usum128[87]),u_counter[5],usum64[43]),u_counter[4],usum32[21]),u_counter[3],usum16[10]),PE(PE(PE(PE(LLR[14],LLR[142],u_counter[6],usum128[88]),PE(LLR[78],LLR[206],u_counter[6],usum128[89]),u_counter[5],usum64[44]),PE(PE(LLR[46],LLR[174],u_counter[6],usum128[90]),PE(LLR[110],LLR[238],u_counter[6],usum128[91]),u_counter[5],usum64[45]),u_counter[4],usum32[22]),PE(PE(PE(LLR[30],LLR[158],u_counter[6],usum128[92]),PE(LLR[94],LLR[222],u_counter[6],usum128[93]),u_counter[5],usum64[46]),PE(PE(LLR[62],LLR[190],u_counter[6],usum128[94]),PE(LLR[126],LLR[254],u_counter[6],usum128[95]),u_counter[5],usum64[47]),u_counter[4],usum32[23]),u_counter[3],usum16[11]),u_counter[2],usum8[5]),u_counter[1],usum4[2]),PE(PE(PE(PE(PE(PE(LLR[4],LLR[132],u_counter[6],usum128[96]),PE(LLR[68],LLR[196],u_counter[6],usum128[97]),u_counter[5],usum64[48]),PE(PE(LLR[36],LLR[164],u_counter[6],usum128[98]),PE(LLR[100],LLR[228],u_counter[6],usum128[99]),u_counter[5],usum64[49]),u_counter[4],usum32[24]),PE(PE(PE(LLR[20],LLR[148],u_counter[6],usum128[100]),PE(LLR[84],LLR[212],u_counter[6],usum128[101]),u_counter[5],usum64[50]),PE(PE(LLR[52],LLR[180],u_counter[6],usum128[102]),PE(LLR[116],LLR[244],u_counter[6],usum128[103]),u_counter[5],usum64[51]),u_counter[4],usum32[25]),u_counter[3],usum16[12]),PE(PE(PE(PE(LLR[12],LLR[140],u_counter[6],usum128[104]),PE(LLR[76],LLR[204],u_counter[6],usum128[105]),u_counter[5],usum64[52]),PE(PE(LLR[44],LLR[172],u_counter[6],usum128[106]),PE(LLR[108],LLR[236],u_counter[6],usum128[107]),u_counter[5],usum64[53]),u_counter[4],usum32[26]),PE(PE(PE(LLR[28],LLR[156],u_counter[6],usum128[108]),PE(LLR[92],LLR[220],u_counter[6],usum128[109]),u_counter[5],usum64[54]),PE(PE(LLR[60],LLR[188],u_counter[6],usum128[110]),PE(LLR[124],LLR[252],u_counter[6],usum128[111]),u_counter[5],usum64[55]),u_counter[4],usum32[27]),u_counter[3],usum16[13]),u_counter[2],usum8[6]),PE(PE(PE(PE(PE(LLR[8],LLR[136],u_counter[6],usum128[112]),PE(LLR[72],LLR[200],u_counter[6],usum128[113]),u_counter[5],usum64[56]),PE(PE(LLR[40],LLR[168],u_counter[6],usum128[114]),PE(LLR[104],LLR[232],u_counter[6],usum128[115]),u_counter[5],usum64[57]),u_counter[4],usum32[28]),PE(PE(PE(LLR[24],LLR[152],u_counter[6],usum128[116]),PE(LLR[88],LLR[216],u_counter[6],usum128[117]),u_counter[5],usum64[58]),PE(PE(LLR[56],LLR[184],u_counter[6],usum128[118]),PE(LLR[120],LLR[248],u_counter[6],usum128[119]),u_counter[5],usum64[59]),u_counter[4],usum32[29]),u_counter[3],usum16[14]),PE(PE(PE(PE(LLR[16],LLR[144],u_counter[6],usum128[120]),PE(LLR[80],LLR[208],u_counter[6],usum128[121]),u_counter[5],usum64[60]),PE(PE(LLR[48],LLR[176],u_counter[6],usum128[122]),PE(LLR[112],LLR[240],u_counter[6],usum128[123]),u_counter[5],usum64[61]),u_counter[4],usum32[30]),PE(PE(PE(LLR[32],LLR[160],u_counter[6],usum128[124]),PE(LLR[96],LLR[224],u_counter[6],usum128[125]),u_counter[5],usum64[62]),PE(PE(LLR[64],LLR[192],u_counter[6],usum128[126]),PE(LLR[128],LLR[256],u_counter[6],usum128[127]),u_counter[5],usum64[63]),u_counter[4],usum32[31]),u_counter[3],usum16[15]),u_counter[2],usum8[7]),u_counter[1],usum4[3]),u_counter[0],usum2[1]);
assign input1_512 = PE(PE(PE(PE(PE(PE(PE(PE(LLR[1],LLR[257],u_counter[7],usum256[0]),PE(LLR[129],LLR[385],u_counter[7],usum256[1]),u_counter[6],usum128[0]),PE(PE(LLR[65],LLR[321],u_counter[7],usum256[2]),PE(LLR[193],LLR[449],u_counter[7],usum256[3]),u_counter[6],usum128[1]),u_counter[5],usum64[0]),PE(PE(PE(LLR[33],LLR[289],u_counter[7],usum256[4]),PE(LLR[161],LLR[417],u_counter[7],usum256[5]),u_counter[6],usum128[2]),PE(PE(LLR[97],LLR[353],u_counter[7],usum256[6]),PE(LLR[225],LLR[481],u_counter[7],usum256[7]),u_counter[6],usum128[3]),u_counter[5],usum64[1]),u_counter[4],usum32[0]),PE(PE(PE(PE(LLR[17],LLR[273],u_counter[7],usum256[8]),PE(LLR[145],LLR[401],u_counter[7],usum256[9]),u_counter[6],usum128[4]),PE(PE(LLR[81],LLR[337],u_counter[7],usum256[10]),PE(LLR[209],LLR[465],u_counter[7],usum256[11]),u_counter[6],usum128[5]),u_counter[5],usum64[2]),PE(PE(PE(LLR[49],LLR[305],u_counter[7],usum256[12]),PE(LLR[177],LLR[433],u_counter[7],usum256[13]),u_counter[6],usum128[6]),PE(PE(LLR[113],LLR[369],u_counter[7],usum256[14]),PE(LLR[241],LLR[497],u_counter[7],usum256[15]),u_counter[6],usum128[7]),u_counter[5],usum64[3]),u_counter[4],usum32[1]),u_counter[3],usum16[0]),PE(PE(PE(PE(PE(LLR[9],LLR[265],u_counter[7],usum256[16]),PE(LLR[137],LLR[393],u_counter[7],usum256[17]),u_counter[6],usum128[8]),PE(PE(LLR[73],LLR[329],u_counter[7],usum256[18]),PE(LLR[201],LLR[457],u_counter[7],usum256[19]),u_counter[6],usum128[9]),u_counter[5],usum64[4]),PE(PE(PE(LLR[41],LLR[297],u_counter[7],usum256[20]),PE(LLR[169],LLR[425],u_counter[7],usum256[21]),u_counter[6],usum128[10]),PE(PE(LLR[105],LLR[361],u_counter[7],usum256[22]),PE(LLR[233],LLR[489],u_counter[7],usum256[23]),u_counter[6],usum128[11]),u_counter[5],usum64[5]),u_counter[4],usum32[2]),PE(PE(PE(PE(LLR[25],LLR[281],u_counter[7],usum256[24]),PE(LLR[153],LLR[409],u_counter[7],usum256[25]),u_counter[6],usum128[12]),PE(PE(LLR[89],LLR[345],u_counter[7],usum256[26]),PE(LLR[217],LLR[473],u_counter[7],usum256[27]),u_counter[6],usum128[13]),u_counter[5],usum64[6]),PE(PE(PE(LLR[57],LLR[313],u_counter[7],usum256[28]),PE(LLR[185],LLR[441],u_counter[7],usum256[29]),u_counter[6],usum128[14]),PE(PE(LLR[121],LLR[377],u_counter[7],usum256[30]),PE(LLR[249],LLR[505],u_counter[7],usum256[31]),u_counter[6],usum128[15]),u_counter[5],usum64[7]),u_counter[4],usum32[3]),u_counter[3],usum16[1]),u_counter[2],usum8[0]),PE(PE(PE(PE(PE(PE(LLR[5],LLR[261],u_counter[7],usum256[32]),PE(LLR[133],LLR[389],u_counter[7],usum256[33]),u_counter[6],usum128[16]),PE(PE(LLR[69],LLR[325],u_counter[7],usum256[34]),PE(LLR[197],LLR[453],u_counter[7],usum256[35]),u_counter[6],usum128[17]),u_counter[5],usum64[8]),PE(PE(PE(LLR[37],LLR[293],u_counter[7],usum256[36]),PE(LLR[165],LLR[421],u_counter[7],usum256[37]),u_counter[6],usum128[18]),PE(PE(LLR[101],LLR[357],u_counter[7],usum256[38]),PE(LLR[229],LLR[485],u_counter[7],usum256[39]),u_counter[6],usum128[19]),u_counter[5],usum64[9]),u_counter[4],usum32[4]),PE(PE(PE(PE(LLR[21],LLR[277],u_counter[7],usum256[40]),PE(LLR[149],LLR[405],u_counter[7],usum256[41]),u_counter[6],usum128[20]),PE(PE(LLR[85],LLR[341],u_counter[7],usum256[42]),PE(LLR[213],LLR[469],u_counter[7],usum256[43]),u_counter[6],usum128[21]),u_counter[5],usum64[10]),PE(PE(PE(LLR[53],LLR[309],u_counter[7],usum256[44]),PE(LLR[181],LLR[437],u_counter[7],usum256[45]),u_counter[6],usum128[22]),PE(PE(LLR[117],LLR[373],u_counter[7],usum256[46]),PE(LLR[245],LLR[501],u_counter[7],usum256[47]),u_counter[6],usum128[23]),u_counter[5],usum64[11]),u_counter[4],usum32[5]),u_counter[3],usum16[2]),PE(PE(PE(PE(PE(LLR[13],LLR[269],u_counter[7],usum256[48]),PE(LLR[141],LLR[397],u_counter[7],usum256[49]),u_counter[6],usum128[24]),PE(PE(LLR[77],LLR[333],u_counter[7],usum256[50]),PE(LLR[205],LLR[461],u_counter[7],usum256[51]),u_counter[6],usum128[25]),u_counter[5],usum64[12]),PE(PE(PE(LLR[45],LLR[301],u_counter[7],usum256[52]),PE(LLR[173],LLR[429],u_counter[7],usum256[53]),u_counter[6],usum128[26]),PE(PE(LLR[109],LLR[365],u_counter[7],usum256[54]),PE(LLR[237],LLR[493],u_counter[7],usum256[55]),u_counter[6],usum128[27]),u_counter[5],usum64[13]),u_counter[4],usum32[6]),PE(PE(PE(PE(LLR[29],LLR[285],u_counter[7],usum256[56]),PE(LLR[157],LLR[413],u_counter[7],usum256[57]),u_counter[6],usum128[28]),PE(PE(LLR[93],LLR[349],u_counter[7],usum256[58]),PE(LLR[221],LLR[477],u_counter[7],usum256[59]),u_counter[6],usum128[29]),u_counter[5],usum64[14]),PE(PE(PE(LLR[61],LLR[317],u_counter[7],usum256[60]),PE(LLR[189],LLR[445],u_counter[7],usum256[61]),u_counter[6],usum128[30]),PE(PE(LLR[125],LLR[381],u_counter[7],usum256[62]),PE(LLR[253],LLR[509],u_counter[7],usum256[63]),u_counter[6],usum128[31]),u_counter[5],usum64[15]),u_counter[4],usum32[7]),u_counter[3],usum16[3]),u_counter[2],usum8[1]),u_counter[1],usum4[0]),PE(PE(PE(PE(PE(PE(PE(LLR[3],LLR[259],u_counter[7],usum256[64]),PE(LLR[131],LLR[387],u_counter[7],usum256[65]),u_counter[6],usum128[32]),PE(PE(LLR[67],LLR[323],u_counter[7],usum256[66]),PE(LLR[195],LLR[451],u_counter[7],usum256[67]),u_counter[6],usum128[33]),u_counter[5],usum64[16]),PE(PE(PE(LLR[35],LLR[291],u_counter[7],usum256[68]),PE(LLR[163],LLR[419],u_counter[7],usum256[69]),u_counter[6],usum128[34]),PE(PE(LLR[99],LLR[355],u_counter[7],usum256[70]),PE(LLR[227],LLR[483],u_counter[7],usum256[71]),u_counter[6],usum128[35]),u_counter[5],usum64[17]),u_counter[4],usum32[8]),PE(PE(PE(PE(LLR[19],LLR[275],u_counter[7],usum256[72]),PE(LLR[147],LLR[403],u_counter[7],usum256[73]),u_counter[6],usum128[36]),PE(PE(LLR[83],LLR[339],u_counter[7],usum256[74]),PE(LLR[211],LLR[467],u_counter[7],usum256[75]),u_counter[6],usum128[37]),u_counter[5],usum64[18]),PE(PE(PE(LLR[51],LLR[307],u_counter[7],usum256[76]),PE(LLR[179],LLR[435],u_counter[7],usum256[77]),u_counter[6],usum128[38]),PE(PE(LLR[115],LLR[371],u_counter[7],usum256[78]),PE(LLR[243],LLR[499],u_counter[7],usum256[79]),u_counter[6],usum128[39]),u_counter[5],usum64[19]),u_counter[4],usum32[9]),u_counter[3],usum16[4]),PE(PE(PE(PE(PE(LLR[11],LLR[267],u_counter[7],usum256[80]),PE(LLR[139],LLR[395],u_counter[7],usum256[81]),u_counter[6],usum128[40]),PE(PE(LLR[75],LLR[331],u_counter[7],usum256[82]),PE(LLR[203],LLR[459],u_counter[7],usum256[83]),u_counter[6],usum128[41]),u_counter[5],usum64[20]),PE(PE(PE(LLR[43],LLR[299],u_counter[7],usum256[84]),PE(LLR[171],LLR[427],u_counter[7],usum256[85]),u_counter[6],usum128[42]),PE(PE(LLR[107],LLR[363],u_counter[7],usum256[86]),PE(LLR[235],LLR[491],u_counter[7],usum256[87]),u_counter[6],usum128[43]),u_counter[5],usum64[21]),u_counter[4],usum32[10]),PE(PE(PE(PE(LLR[27],LLR[283],u_counter[7],usum256[88]),PE(LLR[155],LLR[411],u_counter[7],usum256[89]),u_counter[6],usum128[44]),PE(PE(LLR[91],LLR[347],u_counter[7],usum256[90]),PE(LLR[219],LLR[475],u_counter[7],usum256[91]),u_counter[6],usum128[45]),u_counter[5],usum64[22]),PE(PE(PE(LLR[59],LLR[315],u_counter[7],usum256[92]),PE(LLR[187],LLR[443],u_counter[7],usum256[93]),u_counter[6],usum128[46]),PE(PE(LLR[123],LLR[379],u_counter[7],usum256[94]),PE(LLR[251],LLR[507],u_counter[7],usum256[95]),u_counter[6],usum128[47]),u_counter[5],usum64[23]),u_counter[4],usum32[11]),u_counter[3],usum16[5]),u_counter[2],usum8[2]),PE(PE(PE(PE(PE(PE(LLR[7],LLR[263],u_counter[7],usum256[96]),PE(LLR[135],LLR[391],u_counter[7],usum256[97]),u_counter[6],usum128[48]),PE(PE(LLR[71],LLR[327],u_counter[7],usum256[98]),PE(LLR[199],LLR[455],u_counter[7],usum256[99]),u_counter[6],usum128[49]),u_counter[5],usum64[24]),PE(PE(PE(LLR[39],LLR[295],u_counter[7],usum256[100]),PE(LLR[167],LLR[423],u_counter[7],usum256[101]),u_counter[6],usum128[50]),PE(PE(LLR[103],LLR[359],u_counter[7],usum256[102]),PE(LLR[231],LLR[487],u_counter[7],usum256[103]),u_counter[6],usum128[51]),u_counter[5],usum64[25]),u_counter[4],usum32[12]),PE(PE(PE(PE(LLR[23],LLR[279],u_counter[7],usum256[104]),PE(LLR[151],LLR[407],u_counter[7],usum256[105]),u_counter[6],usum128[52]),PE(PE(LLR[87],LLR[343],u_counter[7],usum256[106]),PE(LLR[215],LLR[471],u_counter[7],usum256[107]),u_counter[6],usum128[53]),u_counter[5],usum64[26]),PE(PE(PE(LLR[55],LLR[311],u_counter[7],usum256[108]),PE(LLR[183],LLR[439],u_counter[7],usum256[109]),u_counter[6],usum128[54]),PE(PE(LLR[119],LLR[375],u_counter[7],usum256[110]),PE(LLR[247],LLR[503],u_counter[7],usum256[111]),u_counter[6],usum128[55]),u_counter[5],usum64[27]),u_counter[4],usum32[13]),u_counter[3],usum16[6]),PE(PE(PE(PE(PE(LLR[15],LLR[271],u_counter[7],usum256[112]),PE(LLR[143],LLR[399],u_counter[7],usum256[113]),u_counter[6],usum128[56]),PE(PE(LLR[79],LLR[335],u_counter[7],usum256[114]),PE(LLR[207],LLR[463],u_counter[7],usum256[115]),u_counter[6],usum128[57]),u_counter[5],usum64[28]),PE(PE(PE(LLR[47],LLR[303],u_counter[7],usum256[116]),PE(LLR[175],LLR[431],u_counter[7],usum256[117]),u_counter[6],usum128[58]),PE(PE(LLR[111],LLR[367],u_counter[7],usum256[118]),PE(LLR[239],LLR[495],u_counter[7],usum256[119]),u_counter[6],usum128[59]),u_counter[5],usum64[29]),u_counter[4],usum32[14]),PE(PE(PE(PE(LLR[31],LLR[287],u_counter[7],usum256[120]),PE(LLR[159],LLR[415],u_counter[7],usum256[121]),u_counter[6],usum128[60]),PE(PE(LLR[95],LLR[351],u_counter[7],usum256[122]),PE(LLR[223],LLR[479],u_counter[7],usum256[123]),u_counter[6],usum128[61]),u_counter[5],usum64[30]),PE(PE(PE(LLR[63],LLR[319],u_counter[7],usum256[124]),PE(LLR[191],LLR[447],u_counter[7],usum256[125]),u_counter[6],usum128[62]),PE(PE(LLR[127],LLR[383],u_counter[7],usum256[126]),PE(LLR[255],LLR[511],u_counter[7],usum256[127]),u_counter[6],usum128[63]),u_counter[5],usum64[31]),u_counter[4],usum32[15]),u_counter[3],usum16[7]),u_counter[2],usum8[3]),u_counter[1],usum4[1]),u_counter[0],usum2[0]);
assign input2_512 = PE(PE(PE(PE(PE(PE(PE(PE(LLR[2],LLR[258],u_counter[7],usum256[128]),PE(LLR[130],LLR[386],u_counter[7],usum256[129]),u_counter[6],usum128[64]),PE(PE(LLR[66],LLR[322],u_counter[7],usum256[130]),PE(LLR[194],LLR[450],u_counter[7],usum256[131]),u_counter[6],usum128[65]),u_counter[5],usum64[32]),PE(PE(PE(LLR[34],LLR[290],u_counter[7],usum256[132]),PE(LLR[162],LLR[418],u_counter[7],usum256[133]),u_counter[6],usum128[66]),PE(PE(LLR[98],LLR[354],u_counter[7],usum256[134]),PE(LLR[226],LLR[482],u_counter[7],usum256[135]),u_counter[6],usum128[67]),u_counter[5],usum64[33]),u_counter[4],usum32[16]),PE(PE(PE(PE(LLR[18],LLR[274],u_counter[7],usum256[136]),PE(LLR[146],LLR[402],u_counter[7],usum256[137]),u_counter[6],usum128[68]),PE(PE(LLR[82],LLR[338],u_counter[7],usum256[138]),PE(LLR[210],LLR[466],u_counter[7],usum256[139]),u_counter[6],usum128[69]),u_counter[5],usum64[34]),PE(PE(PE(LLR[50],LLR[306],u_counter[7],usum256[140]),PE(LLR[178],LLR[434],u_counter[7],usum256[141]),u_counter[6],usum128[70]),PE(PE(LLR[114],LLR[370],u_counter[7],usum256[142]),PE(LLR[242],LLR[498],u_counter[7],usum256[143]),u_counter[6],usum128[71]),u_counter[5],usum64[35]),u_counter[4],usum32[17]),u_counter[3],usum16[8]),PE(PE(PE(PE(PE(LLR[10],LLR[266],u_counter[7],usum256[144]),PE(LLR[138],LLR[394],u_counter[7],usum256[145]),u_counter[6],usum128[72]),PE(PE(LLR[74],LLR[330],u_counter[7],usum256[146]),PE(LLR[202],LLR[458],u_counter[7],usum256[147]),u_counter[6],usum128[73]),u_counter[5],usum64[36]),PE(PE(PE(LLR[42],LLR[298],u_counter[7],usum256[148]),PE(LLR[170],LLR[426],u_counter[7],usum256[149]),u_counter[6],usum128[74]),PE(PE(LLR[106],LLR[362],u_counter[7],usum256[150]),PE(LLR[234],LLR[490],u_counter[7],usum256[151]),u_counter[6],usum128[75]),u_counter[5],usum64[37]),u_counter[4],usum32[18]),PE(PE(PE(PE(LLR[26],LLR[282],u_counter[7],usum256[152]),PE(LLR[154],LLR[410],u_counter[7],usum256[153]),u_counter[6],usum128[76]),PE(PE(LLR[90],LLR[346],u_counter[7],usum256[154]),PE(LLR[218],LLR[474],u_counter[7],usum256[155]),u_counter[6],usum128[77]),u_counter[5],usum64[38]),PE(PE(PE(LLR[58],LLR[314],u_counter[7],usum256[156]),PE(LLR[186],LLR[442],u_counter[7],usum256[157]),u_counter[6],usum128[78]),PE(PE(LLR[122],LLR[378],u_counter[7],usum256[158]),PE(LLR[250],LLR[506],u_counter[7],usum256[159]),u_counter[6],usum128[79]),u_counter[5],usum64[39]),u_counter[4],usum32[19]),u_counter[3],usum16[9]),u_counter[2],usum8[4]),PE(PE(PE(PE(PE(PE(LLR[6],LLR[262],u_counter[7],usum256[160]),PE(LLR[134],LLR[390],u_counter[7],usum256[161]),u_counter[6],usum128[80]),PE(PE(LLR[70],LLR[326],u_counter[7],usum256[162]),PE(LLR[198],LLR[454],u_counter[7],usum256[163]),u_counter[6],usum128[81]),u_counter[5],usum64[40]),PE(PE(PE(LLR[38],LLR[294],u_counter[7],usum256[164]),PE(LLR[166],LLR[422],u_counter[7],usum256[165]),u_counter[6],usum128[82]),PE(PE(LLR[102],LLR[358],u_counter[7],usum256[166]),PE(LLR[230],LLR[486],u_counter[7],usum256[167]),u_counter[6],usum128[83]),u_counter[5],usum64[41]),u_counter[4],usum32[20]),PE(PE(PE(PE(LLR[22],LLR[278],u_counter[7],usum256[168]),PE(LLR[150],LLR[406],u_counter[7],usum256[169]),u_counter[6],usum128[84]),PE(PE(LLR[86],LLR[342],u_counter[7],usum256[170]),PE(LLR[214],LLR[470],u_counter[7],usum256[171]),u_counter[6],usum128[85]),u_counter[5],usum64[42]),PE(PE(PE(LLR[54],LLR[310],u_counter[7],usum256[172]),PE(LLR[182],LLR[438],u_counter[7],usum256[173]),u_counter[6],usum128[86]),PE(PE(LLR[118],LLR[374],u_counter[7],usum256[174]),PE(LLR[246],LLR[502],u_counter[7],usum256[175]),u_counter[6],usum128[87]),u_counter[5],usum64[43]),u_counter[4],usum32[21]),u_counter[3],usum16[10]),PE(PE(PE(PE(PE(LLR[14],LLR[270],u_counter[7],usum256[176]),PE(LLR[142],LLR[398],u_counter[7],usum256[177]),u_counter[6],usum128[88]),PE(PE(LLR[78],LLR[334],u_counter[7],usum256[178]),PE(LLR[206],LLR[462],u_counter[7],usum256[179]),u_counter[6],usum128[89]),u_counter[5],usum64[44]),PE(PE(PE(LLR[46],LLR[302],u_counter[7],usum256[180]),PE(LLR[174],LLR[430],u_counter[7],usum256[181]),u_counter[6],usum128[90]),PE(PE(LLR[110],LLR[366],u_counter[7],usum256[182]),PE(LLR[238],LLR[494],u_counter[7],usum256[183]),u_counter[6],usum128[91]),u_counter[5],usum64[45]),u_counter[4],usum32[22]),PE(PE(PE(PE(LLR[30],LLR[286],u_counter[7],usum256[184]),PE(LLR[158],LLR[414],u_counter[7],usum256[185]),u_counter[6],usum128[92]),PE(PE(LLR[94],LLR[350],u_counter[7],usum256[186]),PE(LLR[222],LLR[478],u_counter[7],usum256[187]),u_counter[6],usum128[93]),u_counter[5],usum64[46]),PE(PE(PE(LLR[62],LLR[318],u_counter[7],usum256[188]),PE(LLR[190],LLR[446],u_counter[7],usum256[189]),u_counter[6],usum128[94]),PE(PE(LLR[126],LLR[382],u_counter[7],usum256[190]),PE(LLR[254],LLR[510],u_counter[7],usum256[191]),u_counter[6],usum128[95]),u_counter[5],usum64[47]),u_counter[4],usum32[23]),u_counter[3],usum16[11]),u_counter[2],usum8[5]),u_counter[1],usum4[2]),PE(PE(PE(PE(PE(PE(PE(LLR[4],LLR[260],u_counter[7],usum256[192]),PE(LLR[132],LLR[388],u_counter[7],usum256[193]),u_counter[6],usum128[96]),PE(PE(LLR[68],LLR[324],u_counter[7],usum256[194]),PE(LLR[196],LLR[452],u_counter[7],usum256[195]),u_counter[6],usum128[97]),u_counter[5],usum64[48]),PE(PE(PE(LLR[36],LLR[292],u_counter[7],usum256[196]),PE(LLR[164],LLR[420],u_counter[7],usum256[197]),u_counter[6],usum128[98]),PE(PE(LLR[100],LLR[356],u_counter[7],usum256[198]),PE(LLR[228],LLR[484],u_counter[7],usum256[199]),u_counter[6],usum128[99]),u_counter[5],usum64[49]),u_counter[4],usum32[24]),PE(PE(PE(PE(LLR[20],LLR[276],u_counter[7],usum256[200]),PE(LLR[148],LLR[404],u_counter[7],usum256[201]),u_counter[6],usum128[100]),PE(PE(LLR[84],LLR[340],u_counter[7],usum256[202]),PE(LLR[212],LLR[468],u_counter[7],usum256[203]),u_counter[6],usum128[101]),u_counter[5],usum64[50]),PE(PE(PE(LLR[52],LLR[308],u_counter[7],usum256[204]),PE(LLR[180],LLR[436],u_counter[7],usum256[205]),u_counter[6],usum128[102]),PE(PE(LLR[116],LLR[372],u_counter[7],usum256[206]),PE(LLR[244],LLR[500],u_counter[7],usum256[207]),u_counter[6],usum128[103]),u_counter[5],usum64[51]),u_counter[4],usum32[25]),u_counter[3],usum16[12]),PE(PE(PE(PE(PE(LLR[12],LLR[268],u_counter[7],usum256[208]),PE(LLR[140],LLR[396],u_counter[7],usum256[209]),u_counter[6],usum128[104]),PE(PE(LLR[76],LLR[332],u_counter[7],usum256[210]),PE(LLR[204],LLR[460],u_counter[7],usum256[211]),u_counter[6],usum128[105]),u_counter[5],usum64[52]),PE(PE(PE(LLR[44],LLR[300],u_counter[7],usum256[212]),PE(LLR[172],LLR[428],u_counter[7],usum256[213]),u_counter[6],usum128[106]),PE(PE(LLR[108],LLR[364],u_counter[7],usum256[214]),PE(LLR[236],LLR[492],u_counter[7],usum256[215]),u_counter[6],usum128[107]),u_counter[5],usum64[53]),u_counter[4],usum32[26]),PE(PE(PE(PE(LLR[28],LLR[284],u_counter[7],usum256[216]),PE(LLR[156],LLR[412],u_counter[7],usum256[217]),u_counter[6],usum128[108]),PE(PE(LLR[92],LLR[348],u_counter[7],usum256[218]),PE(LLR[220],LLR[476],u_counter[7],usum256[219]),u_counter[6],usum128[109]),u_counter[5],usum64[54]),PE(PE(PE(LLR[60],LLR[316],u_counter[7],usum256[220]),PE(LLR[188],LLR[444],u_counter[7],usum256[221]),u_counter[6],usum128[110]),PE(PE(LLR[124],LLR[380],u_counter[7],usum256[222]),PE(LLR[252],LLR[508],u_counter[7],usum256[223]),u_counter[6],usum128[111]),u_counter[5],usum64[55]),u_counter[4],usum32[27]),u_counter[3],usum16[13]),u_counter[2],usum8[6]),PE(PE(PE(PE(PE(PE(LLR[8],LLR[264],u_counter[7],usum256[224]),PE(LLR[136],LLR[392],u_counter[7],usum256[225]),u_counter[6],usum128[112]),PE(PE(LLR[72],LLR[328],u_counter[7],usum256[226]),PE(LLR[200],LLR[456],u_counter[7],usum256[227]),u_counter[6],usum128[113]),u_counter[5],usum64[56]),PE(PE(PE(LLR[40],LLR[296],u_counter[7],usum256[228]),PE(LLR[168],LLR[424],u_counter[7],usum256[229]),u_counter[6],usum128[114]),PE(PE(LLR[104],LLR[360],u_counter[7],usum256[230]),PE(LLR[232],LLR[488],u_counter[7],usum256[231]),u_counter[6],usum128[115]),u_counter[5],usum64[57]),u_counter[4],usum32[28]),PE(PE(PE(PE(LLR[24],LLR[280],u_counter[7],usum256[232]),PE(LLR[152],LLR[408],u_counter[7],usum256[233]),u_counter[6],usum128[116]),PE(PE(LLR[88],LLR[344],u_counter[7],usum256[234]),PE(LLR[216],LLR[472],u_counter[7],usum256[235]),u_counter[6],usum128[117]),u_counter[5],usum64[58]),PE(PE(PE(LLR[56],LLR[312],u_counter[7],usum256[236]),PE(LLR[184],LLR[440],u_counter[7],usum256[237]),u_counter[6],usum128[118]),PE(PE(LLR[120],LLR[376],u_counter[7],usum256[238]),PE(LLR[248],LLR[504],u_counter[7],usum256[239]),u_counter[6],usum128[119]),u_counter[5],usum64[59]),u_counter[4],usum32[29]),u_counter[3],usum16[14]),PE(PE(PE(PE(PE(LLR[16],LLR[272],u_counter[7],usum256[240]),PE(LLR[144],LLR[400],u_counter[7],usum256[241]),u_counter[6],usum128[120]),PE(PE(LLR[80],LLR[336],u_counter[7],usum256[242]),PE(LLR[208],LLR[464],u_counter[7],usum256[243]),u_counter[6],usum128[121]),u_counter[5],usum64[60]),PE(PE(PE(LLR[48],LLR[304],u_counter[7],usum256[244]),PE(LLR[176],LLR[432],u_counter[7],usum256[245]),u_counter[6],usum128[122]),PE(PE(LLR[112],LLR[368],u_counter[7],usum256[246]),PE(LLR[240],LLR[496],u_counter[7],usum256[247]),u_counter[6],usum128[123]),u_counter[5],usum64[61]),u_counter[4],usum32[30]),PE(PE(PE(PE(LLR[32],LLR[288],u_counter[7],usum256[248]),PE(LLR[160],LLR[416],u_counter[7],usum256[249]),u_counter[6],usum128[124]),PE(PE(LLR[96],LLR[352],u_counter[7],usum256[250]),PE(LLR[224],LLR[480],u_counter[7],usum256[251]),u_counter[6],usum128[125]),u_counter[5],usum64[62]),PE(PE(PE(LLR[64],LLR[320],u_counter[7],usum256[252]),PE(LLR[192],LLR[448],u_counter[7],usum256[253]),u_counter[6],usum128[126]),PE(PE(LLR[128],LLR[384],u_counter[7],usum256[254]),PE(LLR[256],LLR[512],u_counter[7],usum256[255]),u_counter[6],usum128[127]),u_counter[5],usum64[63]),u_counter[4],usum32[31]),u_counter[3],usum16[15]),u_counter[2],usum8[7]),u_counter[1],usum4[3]),u_counter[0],usum2[1]);

assign pnode_128 = pnode(input1_128, input2_128, frozen[0], frozen[1]);
assign pnode_256 = pnode(input1_256, input2_256, frozen[0], frozen[1]);
assign pnode_512 = pnode(input1_512, input2_512, frozen[0], frozen[1]);
assign pnode_N   = (N==128) ? pnode_128 : ((N==256) ? pnode_256 : pnode_512);

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		counter_answer <= 0;
		answer <= 0;
	end else if(state==DONE) begin
		counter_answer <= 0;
		answer <= 0;
	end else if(state==DECODE && counter[0]==0 && counter<N) begin
		if(frozen[0] == 0 && frozen[1] == 0) begin
			answer[counter_answer]   <= pnode_N[0];
			answer[counter_answer+1] <= pnode_N[1];
			counter_answer <= counter_answer+2;
		end else if(frozen[0] == 0 && frozen[1] == 1) begin
			answer[counter_answer] <= pnode_N[0];
			counter_answer <= counter_answer+1;
		end else if(frozen[0] == 1 && frozen[1] == 0) begin
			answer[counter_answer] <= pnode_N[1];
			counter_answer <= counter_answer+1;
		end	else begin
			counter_answer <= counter_answer;
		end
	end else begin
		counter_answer <= counter_answer;
		answer <= answer;
	end
end

// **********************//
// *****   OUTPUT   *****//
// **********************//

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		waddr_r     <= 0;
		wdata_r     <= 0;
		proc_done_r <= 0;
	end else if(proc_done_r) begin
		waddr_r     <= 0;
		wdata_r     <= 0;
		proc_done_r <= 0;
	end else begin
		waddr_r     <= (state==DECODE && counter == N-1) ? counter_p : waddr_r;
		wdata_r     <= (state==DECODE && counter == N-1) ? answer : wdata_r;
		proc_done_r <= (!firstRead && state == SUB && counter_p == n_package);
	end
end

assign raddr = (state==SUB) ? 0 :
		       (state==SUB2) ? counter_p*33+counter+1 :
		       (state==READ && counter<=31) ? counter_p*33+counter+2 : 50;
assign waddr = waddr_r;
assign wdata = wdata_r;
assign proc_done = proc_done_r;

// ***********************//
// *****   FUNCTION  *****//
// ***********************//

//***********//
// step1: PE //
//***********//

function [(LLR_bit-2):0] abs;
input signed [(LLR_bit-1):0] x;
abs = (x[(LLR_bit-1)])? -x : x;
endfunction

function [(LLR_bit-1):0] PE;
input [(LLR_bit-1):0] llr_a;
input [(LLR_bit-1):0] llr_b;
input control;
input u_sum;
PE = (control)?	((u_sum) ? (llr_b-llr_a) : (llr_b+llr_a)) :
	 ( llr_a[(LLR_bit-1)]^llr_b[(LLR_bit-1)] ) ?
	 ~( (abs(llr_a)<abs(llr_b))?abs(llr_a):abs(llr_b) )+1 : ( (abs(llr_a)<abs(llr_b))?abs(llr_a):abs(llr_b) );
endfunction

//***************//
// step2: P_NODE //
//***************//

function [1:0] pnode;
input [(LLR_bit-1):0] llr_a;
input [(LLR_bit-1):0] llr_b;
input frozen_a;
input frozen_b;
pnode = {(((llr_b[(LLR_bit-1)] & ~frozen_a) & (((abs(llr_a)>=abs(llr_b))) & ~frozen_b)) |
	   ((((abs(llr_a)>=abs(llr_b))) & ~frozen_b) & (llr_a[(LLR_bit-1)] & frozen_a))) |
	   (llr_b[(LLR_bit-1)] & (~frozen_b & ~((abs(llr_a)>=abs(llr_b))))),
	   (llr_a[(LLR_bit-1)]^llr_b[(LLR_bit-1)]) & ~(frozen_a)};
endfunction

//*******************//
// step3: frozen bit //
//*******************//

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		frozen <= ~(511'b0);
	end else if(state == READ) begin
		frozen[0] <= ( (N==128 && K>=128) ) ? 0 : 1;
		frozen[1] <= ( (N==128 && K>=127) ) ? 0 : 1;
		frozen[2] <= ( (N==128 && K>=126) ) ? 0 : 1;
		frozen[3] <= ( (N==128 && K>=124) ) ? 0 : 1;
		frozen[4] <= ( (N==128 && K>=120) ) ? 0 : 1;
		frozen[5] <= ( (N==128 && K>=112) ) ? 0 : 1;
		frozen[6] <= ( (N==128 && K>=96) ) ? 0 : 1;
		frozen[7] <= ( (N==128 && K>=125) ) ? 0 : 1;
		frozen[8] <= ( (N==128 && K>=123) ) ? 0 : 1;
		frozen[9] <= ( (N==128 && K>=64) ) ? 0 : 1;
		frozen[10] <= ( (N==128 && K>=119) ) ? 0 : 1;
		frozen[11] <= ( (N==128 && K>=122) ) ? 0 : 1;
		frozen[12] <= ( (N==128 && K>=111) ) ? 0 : 1;
		frozen[13] <= ( (N==128 && K>=118) ) ? 0 : 1;
		frozen[14] <= ( (N==128 && K>=110) ) ? 0 : 1;
		frozen[15] <= ( (N==128 && K>=116) || (N==256 && K>=128) ) ? 0 : 1;
		frozen[16] <= ( (N==128 && K>=95) ) ? 0 : 1;
		frozen[17] <= ( (N==128 && K>=63) ) ? 0 : 1;
		frozen[18] <= ( (N==128 && K>=108) ) ? 0 : 1;
		frozen[19] <= ( (N==128 && K>=94) ) ? 0 : 1;
		frozen[20] <= ( (N==128 && K>=104) ) ? 0 : 1;
		frozen[21] <= ( (N==128 && K>=92) ) ? 0 : 1;
		frozen[22] <= ( (N==128 && K>=121) ) ? 0 : 1;
		frozen[23] <= ( (N==128 && K>=62) ) ? 0 : 1;
		frozen[24] <= ( (N==128 && K>=117) || (N==256 && K>=127) ) ? 0 : 1;
		frozen[25] <= ( (N==128 && K>=88) ) ? 0 : 1;
		frozen[26] <= ( (N==128 && K>=60) ) ? 0 : 1;
		frozen[27] <= ( (N==128 && K>=109) ) ? 0 : 1;
		frozen[28] <= ( (N==128 && K>=115) ) ? 0 : 1;
		frozen[29] <= ( (N==128 && K>=80) || (N==256 && K>=126) ) ? 0 : 1;
		frozen[30] <= ( (N==128 && K>=114) ) ? 0 : 1;
		frozen[31] <= ( (N==128 && K>=56) ) ? 0 : 1;
		frozen[32] <= ( (N==128 && K>=107) ) ? 0 : 1;
		frozen[33] <= ( (N==128 && K>=93) ) ? 0 : 1;
		frozen[34] <= ( (N==128 && K>=102) ) ? 0 : 1;
		frozen[35] <= ( (N==128 && K>=48) ) ? 0 : 1;
		frozen[36] <= ( (N==128 && K>=91) || (N==256 && K>=124) ) ? 0 : 1;
		frozen[37] <= ( (N==128 && K>=103) ) ? 0 : 1;
		frozen[38] <= ( (N==128 && K>=106) ) ? 0 : 1;
		frozen[39] <= ( (N==128 && K>=90) ) ? 0 : 1;
		frozen[40] <= ( (N==128 && K>=32) ) ? 0 : 1;
		frozen[41] <= ( (N==128 && K>=61) ) ? 0 : 1;
		frozen[42] <= ( (N==128 && K>=87) ) ? 0 : 1;
		frozen[43] <= ( (N==128 && K>=100) || (N==256 && K>=120) ) ? 0 : 1;
		frozen[44] <= ( (N==128 && K>=59) ) ? 0 : 1;
		frozen[45] <= ( (N==128 && K>=86) ) ? 0 : 1;
		frozen[46] <= ( (N==128 && K>=79) ) ? 0 : 1;
		frozen[47] <= ( (N==128 && K>=54) ) ? 0 : 1;
		frozen[48] <= ( (N==128 && K>=58) || (N==256 && K>=112) ) ? 0 : 1;
		frozen[49] <= ( (N==128 && K>=84) ) ? 0 : 1;
		frozen[50] <= ( (N==128 && K>=47) ) ? 0 : 1;
		frozen[51] <= ( (N==128 && K>=78) ) ? 0 : 1;
		frozen[52] <= ( (N==128 && K>=55) ) ? 0 : 1;
		frozen[53] <= ( (N==128 && K>=113) ) ? 0 : 1;
		frozen[54] <= ( (N==128 && K>=76) || (N==256 && K>=96) ) ? 0 : 1;
		frozen[55] <= ( (N==128 && K>=105) || (N==256 && K>=64) ) ? 0 : 1;
		frozen[56] <= ( (N==128 && K>=52) ) ? 0 : 1;
		frozen[57] <= ( (N==128 && K>=46) ) ? 0 : 1;
		frozen[58] <= ( (N==128 && K>=72) || (N==256 && K>=125) ) ? 0 : 1;
		frozen[59] <= ( (N==128 && K>=101) ) ? 0 : 1;
		frozen[60] <= ( (N==128 && K>=31) ) ? 0 : 1;
		frozen[61] <= ( (N==128 && K>=89) ) ? 0 : 1;
		frozen[62] <= ( (N==128 && K>=44) ) ? 0 : 1;
		frozen[63] <= ( (N==128 && K>=99) || (N==256 && K>=123) ) ? 0 : 1;
		frozen[64] <= ( (N==128 && K>=85) ) ? 0 : 1;
		frozen[65] <= ( (N==128 && K>=30) ) ? 0 : 1;
		frozen[66] <= ( (N==128 && K>=40) || (N==256 && K>=122) ) ? 0 : 1;
		frozen[67] <= ( (N==128 && K>=98) ) ? 0 : 1;
		frozen[68] <= ( (N==128 && K>=57) || (N==256 && K>=119) ) ? 0 : 1;
		frozen[69] <= ( (N==128 && K>=83) ) ? 0 : 1;
		frozen[70] <= ( (N==128 && K>=28) ) ? 0 : 1;
		frozen[71] <= ( (N==128 && K>=77) ) ? 0 : 1;
		frozen[72] <= ( (N==128 && K>=82) ) ? 0 : 1;
		frozen[73] <= ( (N==128 && K>=53) ) ? 0 : 1;
		frozen[74] <= ( (N==128 && K>=24) ) ? 0 : 1;
		frozen[75] <= ( (N==128 && K>=75) || (N==256 && K>=118) || (N==512 && K>=128) ) ? 0 : 1;
		frozen[76] <= ( (N==128 && K>=51) || (N==256 && K>=111) ) ? 0 : 1;
		frozen[77] <= ( (N==128 && K>=74) ) ? 0 : 1;
		frozen[78] <= ( (N==128 && K>=45) ) ? 0 : 1;
		frozen[79] <= ( (N==128 && K>=71) ) ? 0 : 1;
		frozen[80] <= ( (N==128 && K>=16) ) ? 0 : 1;
		frozen[81] <= ( (N==128 && K>=50) || (N==256 && K>=116) ) ? 0 : 1;
		frozen[82] <= ( (N==128 && K>=43) ) ? 0 : 1;
		frozen[83] <= ( (N==128 && K>=70) || (N==256 && K>=110) ) ? 0 : 1;
		frozen[84] <= ( (N==128 && K>=29) ) ? 0 : 1;
		frozen[85] <= ( (N==128 && K>=42) || (N==256 && K>=95) ) ? 0 : 1;
		frozen[86] <= ( (N==128 && K>=68) ) ? 0 : 1;
		frozen[87] <= ( (N==128 && K>=39) ) ? 0 : 1;
		frozen[88] <= ( (N==128 && K>=27) ) ? 0 : 1;
		frozen[89] <= ( (N==128 && K>=97) || (N==256 && K>=108) ) ? 0 : 1;
		frozen[90] <= ( (N==128 && K>=38) ) ? 0 : 1;
		frozen[91] <= ( (N==128 && K>=26) ) ? 0 : 1;
		frozen[92] <= ( (N==128 && K>=23) ) ? 0 : 1;
		frozen[93] <= ( (N==128 && K>=36) || (N==256 && K>=94) ) ? 0 : 1;
		frozen[94] <= ( (N==128 && K>=81) ) ? 0 : 1;
		frozen[95] <= ( (N==128 && K>=22) || (N==256 && K>=63) ) ? 0 : 1;
		frozen[96] <= ( (N==128 && K>=73) || (N==256 && K>=104) ) ? 0 : 1;
		frozen[97] <= ( (N==128 && K>=15) ) ? 0 : 1;
		frozen[98] <= ( (N==128 && K>=49) || (N==256 && K>=92) ) ? 0 : 1;
		frozen[99] <= ( (N==128 && K>=20) ) ? 0 : 1;
		frozen[100] <= ( (N==128 && K>=69) ) ? 0 : 1;
		frozen[101] <= ( (N==128 && K>=14) ) ? 0 : 1;
		frozen[102] <= ( (N==128 && K>=41) ) ? 0 : 1;
		frozen[103] <= ( (N==128 && K>=12) || (N==256 && K>=121) ) ? 0 : 1;
		frozen[104] <= ( (N==128 && K>=67) ) ? 0 : 1;
		frozen[105] <= ( (N==128 && K>=37) || (N==256 && K>=62) ) ? 0 : 1;
		frozen[106] <= ( (N==128 && K>=8) ) ? 0 : 1;
		frozen[107] <= ( (N==128 && K>=66) ) ? 0 : 1;
		frozen[108] <= ( (N==128 && K>=25) || (N==256 && K>=88) ) ? 0 : 1;
		frozen[109] <= ( (N==128 && K>=35) || (N==256 && K>=117) ) ? 0 : 1;
		frozen[110] <= ( (N==128 && K>=21) ) ? 0 : 1;
		frozen[111] <= ( (N==128 && K>=34) ) ? 0 : 1;
		frozen[112] <= ( (N==128 && K>=19) ) ? 0 : 1;
		frozen[113] <= ( (N==128 && K>=13) ) ? 0 : 1;
		frozen[114] <= ( (N==128 && K>=18) || (N==256 && K>=60) ) ? 0 : 1;
		frozen[115] <= ( (N==128 && K>=11) || (N==256 && K>=115) ) ? 0 : 1;
		frozen[116] <= ( (N==128 && K>=10) ) ? 0 : 1;
		frozen[117] <= ( (N==128 && K>=7) || (N==256 && K>=109) ) ? 0 : 1;
		frozen[118] <= ( (N==128 && K>=6) || (N==256 && K>=80) ) ? 0 : 1;
		frozen[119] <= ( (N==128 && K>=65) || (N==256 && K>=114) ) ? 0 : 1;
		frozen[120] <= ( (N==128 && K>=4) ) ? 0 : 1;
		frozen[121] <= ( (N==128 && K>=33) || (N==256 && K>=56) ) ? 0 : 1;
		frozen[122] <= ( (N==128 && K>=17) ) ? 0 : 1;
		frozen[123] <= ( (N==128 && K>=9) || (N==256 && K>=107) ) ? 0 : 1;
		frozen[124] <= ( (N==128 && K>=5) ) ? 0 : 1;
		frozen[125] <= ( (N==128 && K>=3) ) ? 0 : 1;
		frozen[126] <= ( (N==128 && K>=2) || (N==256 && K>=93) ) ? 0 : 1;
		frozen[127] <= ( (N==128 && K>=1) ) ? 0 : 1;
		frozen[128] <= 1;
		frozen[129] <= ( (N==256 && K>=48) ) ? 0 : 1;
		frozen[130] <= ( (N==256 && K>=106) ) ? 0 : 1;
		frozen[131] <= ( (N==256 && K>=103) ) ? 0 : 1;
		frozen[132] <= ( (N==256 && K>=91) ) ? 0 : 1;
		frozen[133] <= 1;
		frozen[134] <= 1;
		frozen[135] <= 1;
		frozen[136] <= ( (N==256 && K>=102) ) ? 0 : 1;
		frozen[137] <= 1;
		frozen[138] <= 1;
		frozen[139] <= ( (N==256 && K>=32) ) ? 0 : 1;
		frozen[140] <= ( (N==256 && K>=90) ) ? 0 : 1;
		frozen[141] <= ( (N==256 && K>=61) ) ? 0 : 1;
		frozen[142] <= 1;
		frozen[143] <= ( (N==256 && K>=87) ) ? 0 : 1;
		frozen[144] <= 1;
		frozen[145] <= ( (N==256 && K>=100) ) ? 0 : 1;
		frozen[146] <= 1;
		frozen[147] <= ( (N==256 && K>=59) ) ? 0 : 1;
		frozen[148] <= ( (N==256 && K>=140) ) ? 0 : 1;
		frozen[149] <= ( (N==256 && K>=86) ) ? 0 : 1;
		frozen[150] <= 1;
		frozen[151] <= ( (N==256 && K>=79) ) ? 0 : 1;
		frozen[152] <= 1;
		frozen[153] <= ( (N==256 && K>=58) ) ? 0 : 1;
		frozen[154] <= ( (N==256 && K>=84) ) ? 0 : 1;
		frozen[155] <= ( (N==256 && K>=136) ) ? 0 : 1;
		frozen[156] <= ( (N==256 && K>=55) ) ? 0 : 1;
		frozen[157] <= ( (N==512 && K>=127) ) ? 0 : 1;
		frozen[158] <= ( (N==256 && K>=113) ) ? 0 : 1;
		frozen[159] <= 1;
		frozen[160] <= ( (N==256 && K>=78) || (N==512 && K>=126) ) ? 0 : 1;
		frozen[161] <= 1;
		frozen[162] <= ( (N==256 && K>=54) ) ? 0 : 1;
		frozen[163] <= 1;
		frozen[164] <= ( (N==256 && K>=76) ) ? 0 : 1;
		frozen[165] <= ( (N==256 && K>=105) ) ? 0 : 1;
		frozen[166] <= ( (N==256 && K>=47) ) ? 0 : 1;
		frozen[167] <= 1;
		frozen[168] <= ( (N==256 && K>=52) ) ? 0 : 1;
		frozen[169] <= ( (N==256 && K>=101) ) ? 0 : 1;
		frozen[170] <= ( (N==256 && K>=46) ) ? 0 : 1;
		frozen[171] <= 1;
		frozen[172] <= ( (N==256 && K>=72) ) ? 0 : 1;
		frozen[173] <= 1;
		frozen[174] <= ( (N==256 && K>=89) ) ? 0 : 1;
		frozen[175] <= ( (N==256 && K>=31) ) ? 0 : 1;
		frozen[176] <= ( (N==256 && K>=99) ) ? 0 : 1;
		frozen[177] <= 1;
		frozen[178] <= ( (N==256 && K>=139) ) ? 0 : 1;
		frozen[179] <= ( (N==256 && K>=44) ) ? 0 : 1;
		frozen[180] <= ( (N==256 && K>=85) ) ? 0 : 1;
		frozen[181] <= ( (N==256 && K>=30) ) ? 0 : 1;
		frozen[182] <= ( (N==256 && K>=40) ) ? 0 : 1;
		frozen[183] <= ( (N==256 && K>=98) ) ? 0 : 1;
		frozen[184] <= ( (N==256 && K>=138) ) ? 0 : 1;
		frozen[185] <= ( (N==256 && K>=83) ) ? 0 : 1;
		frozen[186] <= ( (N==256 && K>=135) ) ? 0 : 1;
		frozen[187] <= ( (N==256 && K>=57) ) ? 0 : 1;
		frozen[188] <= ( (N==256 && K>=77) ) ? 0 : 1;
		frozen[189] <= ( (N==256 && K>=28) ) ? 0 : 1;
		frozen[190] <= ( (N==256 && K>=82) ) ? 0 : 1;
		frozen[191] <= ( (N==256 && K>=134) ) ? 0 : 1;
		frozen[192] <= ( (N==256 && K>=53) || (N==512 && K>=124) ) ? 0 : 1;
		frozen[193] <= 1;
		frozen[194] <= ( (N==256 && K>=75) ) ? 0 : 1;
		frozen[195] <= ( (N==256 && K>=24) ) ? 0 : 1;
		frozen[196] <= ( (N==256 && K>=132) ) ? 0 : 1;
		frozen[197] <= ( (N==256 && K>=51) ) ? 0 : 1;
		frozen[198] <= ( (N==256 && K>=74) ) ? 0 : 1;
		frozen[199] <= ( (N==256 && K>=45) ) ? 0 : 1;
		frozen[200] <= ( (N==256 && K>=71) ) ? 0 : 1;
		frozen[201] <= ( (N==256 && K>=16) ) ? 0 : 1;
		frozen[202] <= ( (N==256 && K>=50) ) ? 0 : 1;
		frozen[203] <= 1;
		frozen[204] <= ( (N==256 && K>=43) ) ? 0 : 1;
		frozen[205] <= ( (N==256 && K>=70) ) ? 0 : 1;
		frozen[206] <= ( (N==256 && K>=29) ) ? 0 : 1;
		frozen[207] <= 1;
		frozen[208] <= ( (N==256 && K>=42) || (N==512 && K>=120) ) ? 0 : 1;
		frozen[209] <= ( (N==256 && K>=68) ) ? 0 : 1;
		frozen[210] <= ( (N==256 && K>=39) ) ? 0 : 1;
		frozen[211] <= ( (N==256 && K>=27) ) ? 0 : 1;
		frozen[212] <= ( (N==256 && K>=97) ) ? 0 : 1;
		frozen[213] <= ( (N==256 && K>=137) ) ? 0 : 1;
		frozen[214] <= ( (N==256 && K>=38) ) ? 0 : 1;
		frozen[215] <= ( (N==256 && K>=26) ) ? 0 : 1;
		frozen[216] <= ( (N==256 && K>=23) ) ? 0 : 1;
		frozen[217] <= ( (N==256 && K>=81) ) ? 0 : 1;
		frozen[218] <= ( (N==256 && K>=133) || (N==512 && K>=112) ) ? 0 : 1;
		frozen[219] <= ( (N==256 && K>=36) ) ? 0 : 1;
		frozen[220] <= ( (N==256 && K>=73) ) ? 0 : 1;
		frozen[221] <= ( (N==256 && K>=22) ) ? 0 : 1;
		frozen[222] <= ( (N==256 && K>=131) ) ? 0 : 1;
		frozen[223] <= ( (N==256 && K>=15) ) ? 0 : 1;
		frozen[224] <= ( (N==256 && K>=49) ) ? 0 : 1;
		frozen[225] <= ( (N==256 && K>=69) ) ? 0 : 1;
		frozen[226] <= ( (N==256 && K>=20) ) ? 0 : 1;
		frozen[227] <= ( (N==256 && K>=130) ) ? 0 : 1;
		frozen[228] <= ( (N==256 && K>=14) ) ? 0 : 1;
		frozen[229] <= ( (N==256 && K>=12) ) ? 0 : 1;
		frozen[230] <= ( (N==256 && K>=67) ) ? 0 : 1;
		frozen[231] <= ( (N==256 && K>=41) ) ? 0 : 1;
		frozen[232] <= ( (N==256 && K>=37) ) ? 0 : 1;
		frozen[233] <= ( (N==256 && K>=25) ) ? 0 : 1;
		frozen[234] <= ( (N==256 && K>=8) ) ? 0 : 1;
		frozen[235] <= ( (N==256 && K>=66) ) ? 0 : 1;
		frozen[236] <= ( (N==256 && K>=35) ) ? 0 : 1;
		frozen[237] <= ( (N==256 && K>=21) ) ? 0 : 1;
		frozen[238] <= ( (N==256 && K>=34) ) ? 0 : 1;
		frozen[239] <= ( (N==256 && K>=19) ) ? 0 : 1;
		frozen[240] <= ( (N==256 && K>=13) || (N==512 && K>=125) ) ? 0 : 1;
		frozen[241] <= ( (N==256 && K>=18) ) ? 0 : 1;
		frozen[242] <= ( (N==256 && K>=11) ) ? 0 : 1;
		frozen[243] <= ( (N==256 && K>=129) || (N==512 && K>=96) ) ? 0 : 1;
		frozen[244] <= ( (N==256 && K>=65) ) ? 0 : 1;
		frozen[245] <= ( (N==256 && K>=10) ) ? 0 : 1;
		frozen[246] <= ( (N==256 && K>=7) ) ? 0 : 1;
		frozen[247] <= ( (N==256 && K>=6) ) ? 0 : 1;
		frozen[248] <= ( (N==256 && K>=4) ) ? 0 : 1;
		frozen[249] <= ( (N==256 && K>=33) ) ? 0 : 1;
		frozen[250] <= ( (N==256 && K>=17) || (N==512 && K>=123) ) ? 0 : 1;
		frozen[251] <= ( (N==256 && K>=5) ) ? 0 : 1;
		frozen[252] <= ( (N==256 && K>=9) ) ? 0 : 1;
		frozen[253] <= ( (N==256 && K>=3) ) ? 0 : 1;
		frozen[254] <= ( (N==256 && K>=2) ) ? 0 : 1;
		frozen[255] <= ( (N==256 && K>=1) ) ? 0 : 1;
		frozen[256] <= 1;
		frozen[257] <= 1;
		frozen[258] <= ( (N==512 && K>=122) ) ? 0 : 1;
		frozen[259] <= 1;
		frozen[260] <= ( (N==512 && K>=119) ) ? 0 : 1;
		frozen[261] <= 1;
		frozen[262] <= 1;
		frozen[263] <= ( (N==512 && K>=64) ) ? 0 : 1;
		frozen[264] <= 1;
		frozen[265] <= 1;
		frozen[266] <= 1;
		frozen[267] <= 1;
		frozen[268] <= ( (N==512 && K>=118) ) ? 0 : 1;
		frozen[269] <= 1;
		frozen[270] <= 1;
		frozen[271] <= 1;
		frozen[272] <= 1;
		frozen[273] <= 1;
		frozen[274] <= 1;
		frozen[275] <= 1;
		frozen[276] <= 1;
		frozen[277] <= 1;
		frozen[278] <= 1;
		frozen[279] <= 1;
		frozen[280] <= ( (N==512 && K>=111) ) ? 0 : 1;
		frozen[281] <= 1;
		frozen[282] <= ( (N==512 && K>=116) ) ? 0 : 1;
		frozen[283] <= 1;
		frozen[284] <= 1;
		frozen[285] <= 1;
		frozen[286] <= 1;
		frozen[287] <= 1;
		frozen[288] <= ( (N==512 && K>=110) ) ? 0 : 1;
		frozen[289] <= 1;
		frozen[290] <= 1;
		frozen[291] <= 1;
		frozen[292] <= ( (N==512 && K>=95) ) ? 0 : 1;
		frozen[293] <= 1;
		frozen[294] <= 1;
		frozen[295] <= ( (N==512 && K>=108) ) ? 0 : 1;
		frozen[296] <= 1;
		frozen[297] <= ( (N==512 && K>=94) ) ? 0 : 1;
		frozen[298] <= 1;
		frozen[299] <= 1;
		frozen[300] <= 1;
		frozen[301] <= 1;
		frozen[302] <= 1;
		frozen[303] <= 1;
		frozen[304] <= 1;
		frozen[305] <= ( (N==512 && K>=63) ) ? 0 : 1;
		frozen[306] <= 1;
		frozen[307] <= ( (N==512 && K>=104) ) ? 0 : 1;
		frozen[308] <= 1;
		frozen[309] <= 1;
		frozen[310] <= ( (N==512 && K>=92) ) ? 0 : 1;
		frozen[311] <= 1;
		frozen[312] <= 1;
		frozen[313] <= 1;
		frozen[314] <= 1;
		frozen[315] <= 1;
		frozen[316] <= 1;
		frozen[317] <= 1;
		frozen[318] <= ( (N==512 && K>=121) ) ? 0 : 1;
		frozen[319] <= 1;
		frozen[320] <= ( (N==512 && K>=62) ) ? 0 : 1;
		frozen[321] <= 1;
		frozen[322] <= 1;
		frozen[323] <= 1;
		frozen[324] <= 1;
		frozen[325] <= 1;
		frozen[326] <= 1;
		frozen[327] <= 1;
		frozen[328] <= ( (N==512 && K>=88) ) ? 0 : 1;
		frozen[329] <= ( (N==512 && K>=117) ) ? 0 : 1;
		frozen[330] <= 1;
		frozen[331] <= 1;
		frozen[332] <= 1;
		frozen[333] <= 1;
		frozen[334] <= 1;
		frozen[335] <= 1;
		frozen[336] <= 1;
		frozen[337] <= 1;
		frozen[338] <= 1;
		frozen[339] <= ( (N==512 && K>=60) ) ? 0 : 1;
		frozen[340] <= ( (N==512 && K>=115) ) ? 0 : 1;
		frozen[341] <= ( (N==512 && K>=109) ) ? 0 : 1;
		frozen[342] <= 1;
		frozen[343] <= ( (N==512 && K>=80) ) ? 0 : 1;
		frozen[344] <= 1;
		frozen[345] <= 1;
		frozen[346] <= 1;
		frozen[347] <= 1;
		frozen[348] <= 1;
		frozen[349] <= ( (N==512 && K>=114) ) ? 0 : 1;
		frozen[350] <= 1;
		frozen[351] <= ( (N==512 && K>=56) ) ? 0 : 1;
		frozen[352] <= 1;
		frozen[353] <= ( (N==512 && K>=107) ) ? 0 : 1;
		frozen[354] <= 1;
		frozen[355] <= 1;
		frozen[356] <= 1;
		frozen[357] <= 1;
		frozen[358] <= 1;
		frozen[359] <= 1;
		frozen[360] <= ( (N==512 && K>=93) ) ? 0 : 1;
		frozen[361] <= ( (N==512 && K>=106) ) ? 0 : 1;
		frozen[362] <= ( (N==512 && K>=48) ) ? 0 : 1;
		frozen[363] <= 1;
		frozen[364] <= ( (N==512 && K>=103) ) ? 0 : 1;
		frozen[365] <= 1;
		frozen[366] <= 1;
		frozen[367] <= ( (N==512 && K>=91) ) ? 0 : 1;
		frozen[368] <= ( (N==512 && K>=102) ) ? 0 : 1;
		frozen[369] <= 1;
		frozen[370] <= 1;
		frozen[371] <= 1;
		frozen[372] <= 1;
		frozen[373] <= 1;
		frozen[374] <= 1;
		frozen[375] <= ( (N==512 && K>=32) ) ? 0 : 1;
		frozen[376] <= 1;
		frozen[377] <= 1;
		frozen[378] <= 1;
		frozen[379] <= ( (N==512 && K>=90) ) ? 0 : 1;
		frozen[380] <= ( (N==512 && K>=87) ) ? 0 : 1;
		frozen[381] <= ( (N==512 && K>=61) ) ? 0 : 1;
		frozen[382] <= 1;
		frozen[383] <= ( (N==512 && K>=100) ) ? 0 : 1;
		frozen[384] <= 1;
		frozen[385] <= ( (N==512 && K>=140) ) ? 0 : 1;
		frozen[386] <= 1;
		frozen[387] <= 1;
		frozen[388] <= ( (N==512 && K>=86) ) ? 0 : 1;
		frozen[389] <= ( (N==512 && K>=59) ) ? 0 : 1;
		frozen[390] <= 1;
		frozen[391] <= ( (N==512 && K>=79) ) ? 0 : 1;
		frozen[392] <= 1;
		frozen[393] <= 1;
		frozen[394] <= ( (N==512 && K>=58) ) ? 0 : 1;
		frozen[395] <= 1;
		frozen[396] <= ( (N==512 && K>=136) ) ? 0 : 1;
		frozen[397] <= ( (N==512 && K>=84) ) ? 0 : 1;
		frozen[398] <= 1;
		frozen[399] <= 1;
		frozen[400] <= ( (N==512 && K>=55) ) ? 0 : 1;
		frozen[401] <= ( (N==512 && K>=113) ) ? 0 : 1;
		frozen[402] <= ( (N==512 && K>=78) ) ? 0 : 1;
		frozen[403] <= 1;
		frozen[404] <= 1;
		frozen[405] <= ( (N==512 && K>=54) ) ? 0 : 1;
		frozen[406] <= 1;
		frozen[407] <= 1;
		frozen[408] <= 1;
		frozen[409] <= ( (N==512 && K>=105) ) ? 0 : 1;
		frozen[410] <= ( (N==512 && K>=76) ) ? 0 : 1;
		frozen[411] <= ( (N==512 && K>=47) ) ? 0 : 1;
		frozen[412] <= 1;
		frozen[413] <= 1;
		frozen[414] <= ( (N==512 && K>=52) ) ? 0 : 1;
		frozen[415] <= 1;
		frozen[416] <= ( (N==512 && K>=101) ) ? 0 : 1;
		frozen[417] <= 1;
		frozen[418] <= ( (N==512 && K>=72) ) ? 0 : 1;
		frozen[419] <= ( (N==512 && K>=138) ) ? 0 : 1;
		frozen[420] <= ( (N==512 && K>=89) ) ? 0 : 1;
		frozen[421] <= ( (N==512 && K>=46) ) ? 0 : 1;
		frozen[422] <= 1;
		frozen[423] <= 1;
		frozen[424] <= ( (N==512 && K>=31) ) ? 0 : 1;
		frozen[425] <= ( (N==512 && K>=99) ) ? 0 : 1;
		frozen[426] <= 1;
		frozen[427] <= ( (N==512 && K>=44) ) ? 0 : 1;
		frozen[428] <= ( (N==512 && K>=83) ) ? 0 : 1;
		frozen[429] <= 1;
		frozen[430] <= ( (N==512 && K>=139) ) ? 0 : 1;
		frozen[431] <= ( (N==512 && K>=30) ) ? 0 : 1;
		frozen[432] <= ( (N==512 && K>=85) ) ? 0 : 1;
		frozen[433] <= ( (N==512 && K>=98) ) ? 0 : 1;
		frozen[434] <= 1;
		frozen[435] <= ( (N==512 && K>=40) ) ? 0 : 1;
		frozen[436] <= ( (N==512 && K>=57) ) ? 0 : 1;
		frozen[437] <= ( (N==512 && K>=135) ) ? 0 : 1;
		frozen[438] <= ( (N==512 && K>=77) ) ? 0 : 1;
		frozen[439] <= 1;
		frozen[440] <= ( (N==512 && K>=28) ) ? 0 : 1;
		frozen[441] <= ( (N==512 && K>=82) ) ? 0 : 1;
		frozen[442] <= ( (N==512 && K>=24) ) ? 0 : 1;
		frozen[443] <= 1;
		frozen[444] <= ( (N==512 && K>=134) ) ? 0 : 1;
		frozen[445] <= ( (N==512 && K>=53) ) ? 0 : 1;
		frozen[446] <= ( (N==512 && K>=75) ) ? 0 : 1;
		frozen[447] <= ( (N==512 && K>=132) ) ? 0 : 1;
		frozen[448] <= ( (N==512 && K>=51) ) ? 0 : 1;
		frozen[449] <= ( (N==512 && K>=16) ) ? 0 : 1;
		frozen[450] <= 1;
		frozen[451] <= ( (N==512 && K>=45) ) ? 0 : 1;
		frozen[452] <= ( (N==512 && K>=74) ) ? 0 : 1;
		frozen[453] <= 1;
		frozen[454] <= ( (N==512 && K>=50) ) ? 0 : 1;
		frozen[455] <= ( (N==512 && K>=70) ) ? 0 : 1;
		frozen[456] <= ( (N==512 && K>=71) ) ? 0 : 1;
		frozen[457] <= ( (N==512 && K>=43) ) ? 0 : 1;
		frozen[458] <= 1;
		frozen[459] <= 1;
		frozen[460] <= 1;
		frozen[461] <= ( (N==512 && K>=137) ) ? 0 : 1;
		frozen[462] <= ( (N==512 && K>=68) ) ? 0 : 1;
		frozen[463] <= ( (N==512 && K>=42) ) ? 0 : 1;
		frozen[464] <= ( (N==512 && K>=29) ) ? 0 : 1;
		frozen[465] <= ( (N==512 && K>=97) ) ? 0 : 1;
		frozen[466] <= ( (N==512 && K>=27) ) ? 0 : 1;
		frozen[467] <= ( (N==512 && K>=39) ) ? 0 : 1;
		frozen[468] <= ( (N==512 && K>=38) ) ? 0 : 1;
		frozen[469] <= 1;
		frozen[470] <= ( (N==512 && K>=133) ) ? 0 : 1;
		frozen[471] <= ( (N==512 && K>=81) ) ? 0 : 1;
		frozen[472] <= ( (N==512 && K>=23) ) ? 0 : 1;
		frozen[473] <= ( (N==512 && K>=26) ) ? 0 : 1;
		frozen[474] <= ( (N==512 && K>=36) ) ? 0 : 1;
		frozen[475] <= ( (N==512 && K>=73) ) ? 0 : 1;
		frozen[476] <= ( (N==512 && K>=22) ) ? 0 : 1;
		frozen[477] <= ( (N==512 && K>=49) ) ? 0 : 1;
		frozen[478] <= ( (N==512 && K>=131) ) ? 0 : 1;
		frozen[479] <= ( (N==512 && K>=15) ) ? 0 : 1;
		frozen[480] <= ( (N==512 && K>=20) ) ? 0 : 1;
		frozen[481] <= ( (N==512 && K>=69) ) ? 0 : 1;
		frozen[482] <= ( (N==512 && K>=130) ) ? 0 : 1;
		frozen[483] <= ( (N==512 && K>=14) ) ? 0 : 1;
		frozen[484] <= ( (N==512 && K>=67) ) ? 0 : 1;
		frozen[485] <= ( (N==512 && K>=41) ) ? 0 : 1;
		frozen[486] <= ( (N==512 && K>=12) ) ? 0 : 1;
		frozen[487] <= ( (N==512 && K>=66) ) ? 0 : 1;
		frozen[488] <= ( (N==512 && K>=37) ) ? 0 : 1;
		frozen[489] <= ( (N==512 && K>=25) ) ? 0 : 1;
		frozen[490] <= ( (N==512 && K>=8) ) ? 0 : 1;
		frozen[491] <= 1;
		frozen[492] <= ( (N==512 && K>=35) ) ? 0 : 1;
		frozen[493] <= ( (N==512 && K>=21) ) ? 0 : 1;
		frozen[494] <= ( (N==512 && K>=34) ) ? 0 : 1;
		frozen[495] <= ( (N==512 && K>=129) ) ? 0 : 1;
		frozen[496] <= ( (N==512 && K>=19) ) ? 0 : 1;
		frozen[497] <= ( (N==512 && K>=13) ) ? 0 : 1;
		frozen[498] <= ( (N==512 && K>=10) ) ? 0 : 1;
		frozen[499] <= ( (N==512 && K>=18) ) ? 0 : 1;
		frozen[500] <= ( (N==512 && K>=11) ) ? 0 : 1;
		frozen[501] <= ( (N==512 && K>=65) ) ? 0 : 1;
		frozen[502] <= ( (N==512 && K>=7) ) ? 0 : 1;
		frozen[503] <= ( (N==512 && K>=6) ) ? 0 : 1;
		frozen[504] <= ( (N==512 && K>=33) ) ? 0 : 1;
		frozen[505] <= ( (N==512 && K>=4) ) ? 0 : 1;
		frozen[506] <= ( (N==512 && K>=17) ) ? 0 : 1;
		frozen[507] <= ( (N==512 && K>=9) ) ? 0 : 1;
		frozen[508] <= ( (N==512 && K>=5) ) ? 0 : 1;
		frozen[509] <= ( (N==512 && K>=3) ) ? 0 : 1;
		frozen[510] <= ( (N==512 && K>=2) ) ? 0 : 1;
		frozen[511] <= ( (N==512 && K>=1) ) ? 0 : 1;
	end else if(state == DECODE && counter[0] == 0 && counter<N) begin
		frozen <= {2'b1,frozen[511:2]};
	end else begin
		frozen <= frozen;
	end
end

endmodule